module Memory(
  input         clock,
  input  [31:0] io_instmem_addr,
  output [31:0] io_instmem_inst,
  input  [31:0] io_datamem_addr,
  output [31:0] io_datamem_rdata,
  input         io_datamem_wen,
  input  [31:0] io_datamem_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [7:0] mem [0:1023]; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_hi_hi_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_instmem_inst_hi_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_hi_lo_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_instmem_inst_hi_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_lo_hi_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_instmem_inst_lo_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_lo_lo_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_instmem_inst_lo_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_hi_hi_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_datamem_rdata_hi_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_hi_lo_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_datamem_rdata_hi_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_lo_hi_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_datamem_rdata_lo_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_lo_lo_data; // @[Memory.scala 45:18]
  wire [9:0] mem_io_datamem_rdata_lo_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_data; // @[Memory.scala 45:18]
  wire [9:0] mem_MPORT_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_1_data; // @[Memory.scala 45:18]
  wire [9:0] mem_MPORT_1_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_1_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_1_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_2_data; // @[Memory.scala 45:18]
  wire [9:0] mem_MPORT_2_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_2_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_2_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_3_data; // @[Memory.scala 45:18]
  wire [9:0] mem_MPORT_3_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_3_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_3_en; // @[Memory.scala 45:18]
  wire [31:0] _io_instmem_inst_T_1 = io_instmem_addr + 32'h3; // @[Memory.scala 51:29]
  wire [31:0] _io_instmem_inst_T_4 = io_instmem_addr + 32'h2; // @[Memory.scala 52:29]
  wire [31:0] _io_instmem_inst_T_7 = io_instmem_addr + 32'h1; // @[Memory.scala 53:29]
  wire [15:0] io_instmem_inst_lo = {mem_io_instmem_inst_lo_hi_data,mem_io_instmem_inst_lo_lo_data}; // @[Cat.scala 30:58]
  wire [15:0] io_instmem_inst_hi = {mem_io_instmem_inst_hi_hi_data,mem_io_instmem_inst_hi_lo_data}; // @[Cat.scala 30:58]
  wire [31:0] _io_datamem_rdata_T_1 = io_datamem_addr + 32'h3; // @[Memory.scala 58:29]
  wire [31:0] _io_datamem_rdata_T_4 = io_datamem_addr + 32'h2; // @[Memory.scala 59:29]
  wire [31:0] _io_datamem_rdata_T_7 = io_datamem_addr + 32'h1; // @[Memory.scala 60:29]
  wire [15:0] io_datamem_rdata_lo = {mem_io_datamem_rdata_lo_hi_data,mem_io_datamem_rdata_lo_lo_data}; // @[Cat.scala 30:58]
  wire [15:0] io_datamem_rdata_hi = {mem_io_datamem_rdata_hi_hi_data,mem_io_datamem_rdata_hi_lo_data}; // @[Cat.scala 30:58]
  assign mem_io_instmem_inst_hi_hi_addr = _io_instmem_inst_T_1[9:0];
  assign mem_io_instmem_inst_hi_hi_data = mem[mem_io_instmem_inst_hi_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_hi_lo_addr = _io_instmem_inst_T_4[9:0];
  assign mem_io_instmem_inst_hi_lo_data = mem[mem_io_instmem_inst_hi_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_lo_hi_addr = _io_instmem_inst_T_7[9:0];
  assign mem_io_instmem_inst_lo_hi_data = mem[mem_io_instmem_inst_lo_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_lo_lo_addr = io_instmem_addr[9:0];
  assign mem_io_instmem_inst_lo_lo_data = mem[mem_io_instmem_inst_lo_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_hi_hi_addr = _io_datamem_rdata_T_1[9:0];
  assign mem_io_datamem_rdata_hi_hi_data = mem[mem_io_datamem_rdata_hi_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_hi_lo_addr = _io_datamem_rdata_T_4[9:0];
  assign mem_io_datamem_rdata_hi_lo_data = mem[mem_io_datamem_rdata_hi_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_lo_hi_addr = _io_datamem_rdata_T_7[9:0];
  assign mem_io_datamem_rdata_lo_hi_data = mem[mem_io_datamem_rdata_lo_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_lo_lo_addr = io_datamem_addr[9:0];
  assign mem_io_datamem_rdata_lo_lo_data = mem[mem_io_datamem_rdata_lo_lo_addr]; // @[Memory.scala 45:18]
  assign mem_MPORT_data = io_datamem_wdata[7:0];
  assign mem_MPORT_addr = io_datamem_addr[9:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_datamem_wen;
  assign mem_MPORT_1_data = io_datamem_wdata[15:8];
  assign mem_MPORT_1_addr = _io_datamem_rdata_T_7[9:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = io_datamem_wen;
  assign mem_MPORT_2_data = io_datamem_wdata[23:16];
  assign mem_MPORT_2_addr = _io_datamem_rdata_T_4[9:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = io_datamem_wen;
  assign mem_MPORT_3_data = io_datamem_wdata[31:24];
  assign mem_MPORT_3_addr = _io_datamem_rdata_T_1[9:0];
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = io_datamem_wen;
  assign io_instmem_inst = {io_instmem_inst_hi,io_instmem_inst_lo}; // @[Cat.scala 30:58]
  assign io_datamem_rdata = {io_datamem_rdata_hi,io_datamem_rdata_lo}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[Memory.scala 45:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PC(
  input         clock,
  input         reset,
  input         io_in_stall_in_stall_flag,
  input  [31:0] io_in_ex_in_alu_out,
  input         io_in_ex_in_jump_flag,
  input         io_in_br_in_br_flag,
  input  [31:0] io_in_br_in_br_target,
  output [31:0] io_out_reg_pc,
  output [31:0] io_out_inst,
  output        io_out_br_flag,
  output        io_out_jump_flag,
  output [31:0] io_instmem_addr,
  input  [31:0] io_instmem_inst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PC.scala 100:38]
  wire [31:0] reg_pc_next_default = reg_pc + 32'h4; // @[PC.scala 101:38]
  wire  _T_1 = ~reset; // @[PC.scala 118:11]
  assign io_out_reg_pc = reg_pc; // @[PC.scala 112:25]
  assign io_out_inst = io_instmem_inst; // @[PC.scala 113:25]
  assign io_out_br_flag = io_in_br_in_br_flag; // @[PC.scala 114:25]
  assign io_out_jump_flag = io_in_ex_in_jump_flag; // @[PC.scala 115:25]
  assign io_instmem_addr = reg_pc; // @[PC.scala 111:25]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 100:38]
      reg_pc <= 32'h0; // @[PC.scala 100:38]
    end else if (io_in_br_in_br_flag) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_br_in_br_target;
    end else if (io_in_ex_in_jump_flag) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_ex_in_alu_out;
    end else if (!(io_in_stall_in_stall_flag)) begin // @[Mux.scala 98:16]
      reg_pc <= reg_pc_next_default;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-----------------------START----------------------\n"); // @[PC.scala 118:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"-------------IF------------\n"); // @[PC.scala 119:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"reg_pc: 0x%x\n",reg_pc); // @[PC.scala 120:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"inst: 0x%x\n",io_instmem_inst); // @[PC.scala 121:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ID(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_in_reg_pc,
  input  [31:0] io_in_if_in_inst,
  input         io_in_if_in_br_flag,
  input         io_in_if_in_jump_flag,
  input         io_in_stall_in_stall_flag,
  input         io_in_mem_in_rd_wen,
  input  [4:0]  io_in_mem_in_rd_addr,
  input  [31:0] io_in_mem_in_rd_data,
  input         io_in_wb_in_rd_wen,
  input  [4:0]  io_in_wb_in_rd_addr,
  input  [31:0] io_in_wb_in_rd_data,
  output [31:0] io_out_op1_data,
  output [31:0] io_out_op2_data,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_csr_addr_default,
  output [4:0]  io_out_exe_fun,
  output        io_out_mem_wen,
  output        io_out_rd_wen,
  output [2:0]  io_out_rd_sel,
  output [2:0]  io_out_csr_cmd,
  output [31:0] io_out_rs2_data,
  output [31:0] io_out_imm_b_sext
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_x_0; // @[ID.scala 75:26]
  reg [31:0] reg_x_1; // @[ID.scala 75:26]
  reg [31:0] reg_x_2; // @[ID.scala 75:26]
  reg [31:0] reg_x_3; // @[ID.scala 75:26]
  reg [31:0] reg_x_4; // @[ID.scala 75:26]
  reg [31:0] reg_x_5; // @[ID.scala 75:26]
  reg [31:0] reg_x_6; // @[ID.scala 75:26]
  reg [31:0] reg_x_7; // @[ID.scala 75:26]
  reg [31:0] reg_x_8; // @[ID.scala 75:26]
  reg [31:0] reg_x_9; // @[ID.scala 75:26]
  reg [31:0] reg_x_10; // @[ID.scala 75:26]
  reg [31:0] reg_x_11; // @[ID.scala 75:26]
  reg [31:0] reg_x_12; // @[ID.scala 75:26]
  reg [31:0] reg_x_13; // @[ID.scala 75:26]
  reg [31:0] reg_x_14; // @[ID.scala 75:26]
  reg [31:0] reg_x_15; // @[ID.scala 75:26]
  reg [31:0] reg_x_16; // @[ID.scala 75:26]
  reg [31:0] reg_x_17; // @[ID.scala 75:26]
  reg [31:0] reg_x_18; // @[ID.scala 75:26]
  reg [31:0] reg_x_19; // @[ID.scala 75:26]
  reg [31:0] reg_x_20; // @[ID.scala 75:26]
  reg [31:0] reg_x_21; // @[ID.scala 75:26]
  reg [31:0] reg_x_22; // @[ID.scala 75:26]
  reg [31:0] reg_x_23; // @[ID.scala 75:26]
  reg [31:0] reg_x_24; // @[ID.scala 75:26]
  reg [31:0] reg_x_25; // @[ID.scala 75:26]
  reg [31:0] reg_x_26; // @[ID.scala 75:26]
  reg [31:0] reg_x_27; // @[ID.scala 75:26]
  reg [31:0] reg_x_28; // @[ID.scala 75:26]
  reg [31:0] reg_x_29; // @[ID.scala 75:26]
  reg [31:0] reg_x_30; // @[ID.scala 75:26]
  reg [31:0] reg_x_31; // @[ID.scala 75:26]
  wire  _inst_T_1 = io_in_if_in_br_flag | io_in_if_in_jump_flag | io_in_stall_in_stall_flag; // @[ID.scala 91:31]
  wire [31:0] inst = _inst_T_1 ? 32'h13 : io_in_if_in_inst; // @[Mux.scala 98:16]
  wire [4:0] rs1_addr = inst[19:15]; // @[ID.scala 95:24]
  wire [4:0] rs2_addr = inst[24:20]; // @[ID.scala 96:24]
  wire [4:0] rd_addr = inst[11:7]; // @[ID.scala 97:24]
  wire [11:0] csr_addr_default = inst[31:20]; // @[ID.scala 98:32]
  wire  _rs1_data_T = rs1_addr == 5'h0; // @[ID.scala 100:19]
  wire  _rs1_data_T_3 = rs1_addr == io_in_mem_in_rd_addr & io_in_mem_in_rd_wen; // @[ID.scala 101:37]
  wire  _rs1_data_T_6 = rs1_addr == io_in_wb_in_rd_addr & io_in_wb_in_rd_wen; // @[ID.scala 102:36]
  wire [31:0] _GEN_1 = 5'h1 == rs1_addr ? reg_x_1 : reg_x_0; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_2 = 5'h2 == rs1_addr ? reg_x_2 : _GEN_1; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_3 = 5'h3 == rs1_addr ? reg_x_3 : _GEN_2; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_4 = 5'h4 == rs1_addr ? reg_x_4 : _GEN_3; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_5 = 5'h5 == rs1_addr ? reg_x_5 : _GEN_4; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_6 = 5'h6 == rs1_addr ? reg_x_6 : _GEN_5; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_7 = 5'h7 == rs1_addr ? reg_x_7 : _GEN_6; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_8 = 5'h8 == rs1_addr ? reg_x_8 : _GEN_7; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_9 = 5'h9 == rs1_addr ? reg_x_9 : _GEN_8; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_10 = 5'ha == rs1_addr ? reg_x_10 : _GEN_9; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_11 = 5'hb == rs1_addr ? reg_x_11 : _GEN_10; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_12 = 5'hc == rs1_addr ? reg_x_12 : _GEN_11; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_13 = 5'hd == rs1_addr ? reg_x_13 : _GEN_12; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_14 = 5'he == rs1_addr ? reg_x_14 : _GEN_13; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_15 = 5'hf == rs1_addr ? reg_x_15 : _GEN_14; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_16 = 5'h10 == rs1_addr ? reg_x_16 : _GEN_15; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_17 = 5'h11 == rs1_addr ? reg_x_17 : _GEN_16; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_18 = 5'h12 == rs1_addr ? reg_x_18 : _GEN_17; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_19 = 5'h13 == rs1_addr ? reg_x_19 : _GEN_18; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_20 = 5'h14 == rs1_addr ? reg_x_20 : _GEN_19; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_21 = 5'h15 == rs1_addr ? reg_x_21 : _GEN_20; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_22 = 5'h16 == rs1_addr ? reg_x_22 : _GEN_21; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_23 = 5'h17 == rs1_addr ? reg_x_23 : _GEN_22; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_24 = 5'h18 == rs1_addr ? reg_x_24 : _GEN_23; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_25 = 5'h19 == rs1_addr ? reg_x_25 : _GEN_24; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_26 = 5'h1a == rs1_addr ? reg_x_26 : _GEN_25; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_27 = 5'h1b == rs1_addr ? reg_x_27 : _GEN_26; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_28 = 5'h1c == rs1_addr ? reg_x_28 : _GEN_27; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_29 = 5'h1d == rs1_addr ? reg_x_29 : _GEN_28; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_30 = 5'h1e == rs1_addr ? reg_x_30 : _GEN_29; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_31 = 5'h1f == rs1_addr ? reg_x_31 : _GEN_30; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _rs1_data_T_7 = _rs1_data_T_6 ? io_in_wb_in_rd_data : _GEN_31; // @[Mux.scala 98:16]
  wire [31:0] _rs1_data_T_8 = _rs1_data_T_3 ? io_in_mem_in_rd_data : _rs1_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] rs1_data = _rs1_data_T ? 32'h0 : _rs1_data_T_8; // @[Mux.scala 98:16]
  wire  _rs2_data_T = rs2_addr == 5'h0; // @[ID.scala 105:19]
  wire  _rs2_data_T_3 = rs2_addr == io_in_mem_in_rd_addr & io_in_mem_in_rd_wen; // @[ID.scala 106:37]
  wire  _rs2_data_T_6 = rs2_addr == io_in_wb_in_rd_addr & io_in_wb_in_rd_wen; // @[ID.scala 107:36]
  wire [31:0] _GEN_33 = 5'h1 == rs2_addr ? reg_x_1 : reg_x_0; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_34 = 5'h2 == rs2_addr ? reg_x_2 : _GEN_33; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_35 = 5'h3 == rs2_addr ? reg_x_3 : _GEN_34; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_36 = 5'h4 == rs2_addr ? reg_x_4 : _GEN_35; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_37 = 5'h5 == rs2_addr ? reg_x_5 : _GEN_36; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_38 = 5'h6 == rs2_addr ? reg_x_6 : _GEN_37; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_39 = 5'h7 == rs2_addr ? reg_x_7 : _GEN_38; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_40 = 5'h8 == rs2_addr ? reg_x_8 : _GEN_39; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_41 = 5'h9 == rs2_addr ? reg_x_9 : _GEN_40; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_42 = 5'ha == rs2_addr ? reg_x_10 : _GEN_41; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_43 = 5'hb == rs2_addr ? reg_x_11 : _GEN_42; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_44 = 5'hc == rs2_addr ? reg_x_12 : _GEN_43; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_45 = 5'hd == rs2_addr ? reg_x_13 : _GEN_44; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_46 = 5'he == rs2_addr ? reg_x_14 : _GEN_45; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_47 = 5'hf == rs2_addr ? reg_x_15 : _GEN_46; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_48 = 5'h10 == rs2_addr ? reg_x_16 : _GEN_47; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_49 = 5'h11 == rs2_addr ? reg_x_17 : _GEN_48; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_50 = 5'h12 == rs2_addr ? reg_x_18 : _GEN_49; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_51 = 5'h13 == rs2_addr ? reg_x_19 : _GEN_50; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_52 = 5'h14 == rs2_addr ? reg_x_20 : _GEN_51; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_53 = 5'h15 == rs2_addr ? reg_x_21 : _GEN_52; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_54 = 5'h16 == rs2_addr ? reg_x_22 : _GEN_53; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_55 = 5'h17 == rs2_addr ? reg_x_23 : _GEN_54; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_56 = 5'h18 == rs2_addr ? reg_x_24 : _GEN_55; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_57 = 5'h19 == rs2_addr ? reg_x_25 : _GEN_56; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_58 = 5'h1a == rs2_addr ? reg_x_26 : _GEN_57; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_59 = 5'h1b == rs2_addr ? reg_x_27 : _GEN_58; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_60 = 5'h1c == rs2_addr ? reg_x_28 : _GEN_59; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_61 = 5'h1d == rs2_addr ? reg_x_29 : _GEN_60; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_62 = 5'h1e == rs2_addr ? reg_x_30 : _GEN_61; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_63 = 5'h1f == rs2_addr ? reg_x_31 : _GEN_62; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _rs2_data_T_7 = _rs2_data_T_6 ? io_in_wb_in_rd_data : _GEN_63; // @[Mux.scala 98:16]
  wire [31:0] _rs2_data_T_8 = _rs2_data_T_3 ? io_in_mem_in_rd_data : _rs2_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] rs2_data = _rs2_data_T ? 32'h0 : _rs2_data_T_8; // @[Mux.scala 98:16]
  wire [19:0] imm_i_sext_hi = csr_addr_default[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_i_sext = {imm_i_sext_hi,csr_addr_default}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi = inst[31:25]; // @[ID.scala 111:31]
  wire [11:0] imm_s = {imm_s_hi,rd_addr}; // @[Cat.scala 30:58]
  wire [19:0] imm_s_sext_hi = imm_s[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_s_sext = {imm_s_sext_hi,imm_s_hi,rd_addr}; // @[Cat.scala 30:58]
  wire  imm_b_hi_hi = inst[31]; // @[ID.scala 113:31]
  wire  imm_b_hi_lo = inst[7]; // @[ID.scala 113:41]
  wire [5:0] imm_b_lo_hi = inst[30:25]; // @[ID.scala 113:50]
  wire [3:0] imm_b_lo_lo = inst[11:8]; // @[ID.scala 113:64]
  wire [11:0] imm_b = {imm_b_hi_hi,imm_b_hi_lo,imm_b_lo_hi,imm_b_lo_lo}; // @[Cat.scala 30:58]
  wire [18:0] imm_b_sext_hi_hi = imm_b[11] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [30:0] imm_b_sext_hi = {imm_b_sext_hi_hi,imm_b_hi_hi,imm_b_hi_lo,imm_b_lo_hi,imm_b_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] imm_j_hi_lo = inst[19:12]; // @[ID.scala 115:41]
  wire  imm_j_lo_hi = inst[20]; // @[ID.scala 115:55]
  wire [9:0] imm_j_lo_lo = inst[30:21]; // @[ID.scala 115:65]
  wire [19:0] imm_j = {imm_b_hi_hi,imm_j_hi_lo,imm_j_lo_hi,imm_j_lo_lo}; // @[Cat.scala 30:58]
  wire [10:0] imm_j_sext_hi_hi = imm_j[19] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_j_sext = {imm_j_sext_hi_hi,imm_b_hi_hi,imm_j_hi_lo,imm_j_lo_hi,imm_j_lo_lo,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] imm_u = inst[31:12]; // @[ID.scala 117:27]
  wire [31:0] imm_u_shifted = {imm_u,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_z_uext = {27'h0,rs1_addr}; // @[Cat.scala 30:58]
  wire [31:0] _inst_type_T = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_4 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h33 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h40000033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h7033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h6033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h4033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h1033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h5033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h40005033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h1013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h5013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h40005013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h2033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h3033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_54 = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h6f == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h37 == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h17 == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h5073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h6073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h7073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire [4:0] _inst_type_T_77 = _inst_type_T_73 ? 5'h12 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_78 = _inst_type_T_71 ? 5'h12 : _inst_type_T_77; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_79 = _inst_type_T_69 ? 5'h12 : _inst_type_T_78; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_80 = _inst_type_T_67 ? 5'h12 : _inst_type_T_79; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_81 = _inst_type_T_65 ? 5'h12 : _inst_type_T_80; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_82 = _inst_type_T_63 ? 5'h12 : _inst_type_T_81; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_83 = _inst_type_T_61 ? 5'h1 : _inst_type_T_82; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_84 = _inst_type_T_59 ? 5'h1 : _inst_type_T_83; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_85 = _inst_type_T_57 ? 5'h11 : _inst_type_T_84; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_86 = _inst_type_T_55 ? 5'h1 : _inst_type_T_85; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_87 = _inst_type_T_53 ? 5'hf : _inst_type_T_86; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_88 = _inst_type_T_51 ? 5'hd : _inst_type_T_87; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_89 = _inst_type_T_49 ? 5'h10 : _inst_type_T_88; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_90 = _inst_type_T_47 ? 5'he : _inst_type_T_89; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_91 = _inst_type_T_45 ? 5'hc : _inst_type_T_90; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_92 = _inst_type_T_43 ? 5'hb : _inst_type_T_91; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_93 = _inst_type_T_41 ? 5'ha : _inst_type_T_92; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_94 = _inst_type_T_39 ? 5'h9 : _inst_type_T_93; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_95 = _inst_type_T_37 ? 5'ha : _inst_type_T_94; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_96 = _inst_type_T_35 ? 5'h9 : _inst_type_T_95; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_97 = _inst_type_T_33 ? 5'h8 : _inst_type_T_96; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_98 = _inst_type_T_31 ? 5'h7 : _inst_type_T_97; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_99 = _inst_type_T_29 ? 5'h6 : _inst_type_T_98; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_100 = _inst_type_T_27 ? 5'h8 : _inst_type_T_99; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_101 = _inst_type_T_25 ? 5'h7 : _inst_type_T_100; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_102 = _inst_type_T_23 ? 5'h6 : _inst_type_T_101; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_103 = _inst_type_T_21 ? 5'h5 : _inst_type_T_102; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_104 = _inst_type_T_19 ? 5'h4 : _inst_type_T_103; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_105 = _inst_type_T_17 ? 5'h3 : _inst_type_T_104; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_106 = _inst_type_T_15 ? 5'h5 : _inst_type_T_105; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_107 = _inst_type_T_13 ? 5'h4 : _inst_type_T_106; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_108 = _inst_type_T_11 ? 5'h3 : _inst_type_T_107; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_109 = _inst_type_T_9 ? 5'h2 : _inst_type_T_108; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_110 = _inst_type_T_7 ? 5'h1 : _inst_type_T_109; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_111 = _inst_type_T_5 ? 5'h1 : _inst_type_T_110; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_112 = _inst_type_T_3 ? 5'h1 : _inst_type_T_111; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_113 = _inst_type_T_75 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_114 = _inst_type_T_73 ? 2'h3 : _inst_type_T_113; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_115 = _inst_type_T_71 ? 2'h0 : _inst_type_T_114; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_116 = _inst_type_T_69 ? 2'h3 : _inst_type_T_115; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_117 = _inst_type_T_67 ? 2'h0 : _inst_type_T_116; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_118 = _inst_type_T_65 ? 2'h3 : _inst_type_T_117; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_119 = _inst_type_T_63 ? 2'h0 : _inst_type_T_118; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_120 = _inst_type_T_61 ? 2'h1 : _inst_type_T_119; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_121 = _inst_type_T_59 ? 2'h2 : _inst_type_T_120; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_122 = _inst_type_T_57 ? 2'h0 : _inst_type_T_121; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_123 = _inst_type_T_55 ? 2'h1 : _inst_type_T_122; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_124 = _inst_type_T_53 ? 2'h0 : _inst_type_T_123; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_125 = _inst_type_T_51 ? 2'h0 : _inst_type_T_124; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_126 = _inst_type_T_49 ? 2'h0 : _inst_type_T_125; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_127 = _inst_type_T_47 ? 2'h0 : _inst_type_T_126; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_128 = _inst_type_T_45 ? 2'h0 : _inst_type_T_127; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_129 = _inst_type_T_43 ? 2'h0 : _inst_type_T_128; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_130 = _inst_type_T_41 ? 2'h0 : _inst_type_T_129; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_131 = _inst_type_T_39 ? 2'h0 : _inst_type_T_130; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_132 = _inst_type_T_37 ? 2'h0 : _inst_type_T_131; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_133 = _inst_type_T_35 ? 2'h0 : _inst_type_T_132; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_134 = _inst_type_T_33 ? 2'h0 : _inst_type_T_133; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_135 = _inst_type_T_31 ? 2'h0 : _inst_type_T_134; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_136 = _inst_type_T_29 ? 2'h0 : _inst_type_T_135; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_137 = _inst_type_T_27 ? 2'h0 : _inst_type_T_136; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_138 = _inst_type_T_25 ? 2'h0 : _inst_type_T_137; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_139 = _inst_type_T_23 ? 2'h0 : _inst_type_T_138; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_140 = _inst_type_T_21 ? 2'h0 : _inst_type_T_139; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_141 = _inst_type_T_19 ? 2'h0 : _inst_type_T_140; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_142 = _inst_type_T_17 ? 2'h0 : _inst_type_T_141; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_143 = _inst_type_T_15 ? 2'h0 : _inst_type_T_142; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_144 = _inst_type_T_13 ? 2'h0 : _inst_type_T_143; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_145 = _inst_type_T_11 ? 2'h0 : _inst_type_T_144; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_146 = _inst_type_T_9 ? 2'h0 : _inst_type_T_145; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_147 = _inst_type_T_7 ? 2'h0 : _inst_type_T_146; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_148 = _inst_type_T_5 ? 2'h0 : _inst_type_T_147; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_149 = _inst_type_T_3 ? 2'h0 : _inst_type_T_148; // @[Lookup.scala 33:37]
  wire [1:0] inst_type_1 = _inst_type_T_1 ? 2'h0 : _inst_type_T_149; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_150 = _inst_type_T_75 ? 3'h0 : 3'h1; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_151 = _inst_type_T_73 ? 3'h0 : _inst_type_T_150; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_152 = _inst_type_T_71 ? 3'h0 : _inst_type_T_151; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_153 = _inst_type_T_69 ? 3'h0 : _inst_type_T_152; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_154 = _inst_type_T_67 ? 3'h0 : _inst_type_T_153; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_155 = _inst_type_T_65 ? 3'h0 : _inst_type_T_154; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_156 = _inst_type_T_63 ? 3'h0 : _inst_type_T_155; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_157 = _inst_type_T_61 ? 3'h5 : _inst_type_T_156; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_158 = _inst_type_T_59 ? 3'h5 : _inst_type_T_157; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_159 = _inst_type_T_57 ? 3'h2 : _inst_type_T_158; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_160 = _inst_type_T_55 ? 3'h4 : _inst_type_T_159; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_161 = _inst_type_T_53 ? 3'h1 : _inst_type_T_160; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_162 = _inst_type_T_51 ? 3'h1 : _inst_type_T_161; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_163 = _inst_type_T_49 ? 3'h1 : _inst_type_T_162; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_164 = _inst_type_T_47 ? 3'h1 : _inst_type_T_163; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_165 = _inst_type_T_45 ? 3'h1 : _inst_type_T_164; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_166 = _inst_type_T_43 ? 3'h1 : _inst_type_T_165; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_167 = _inst_type_T_41 ? 3'h2 : _inst_type_T_166; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_168 = _inst_type_T_39 ? 3'h2 : _inst_type_T_167; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_169 = _inst_type_T_37 ? 3'h1 : _inst_type_T_168; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_170 = _inst_type_T_35 ? 3'h1 : _inst_type_T_169; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_171 = _inst_type_T_33 ? 3'h2 : _inst_type_T_170; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_172 = _inst_type_T_31 ? 3'h2 : _inst_type_T_171; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_173 = _inst_type_T_29 ? 3'h2 : _inst_type_T_172; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_174 = _inst_type_T_27 ? 3'h1 : _inst_type_T_173; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_175 = _inst_type_T_25 ? 3'h1 : _inst_type_T_174; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_176 = _inst_type_T_23 ? 3'h1 : _inst_type_T_175; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_177 = _inst_type_T_21 ? 3'h2 : _inst_type_T_176; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_178 = _inst_type_T_19 ? 3'h2 : _inst_type_T_177; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_179 = _inst_type_T_17 ? 3'h2 : _inst_type_T_178; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_180 = _inst_type_T_15 ? 3'h1 : _inst_type_T_179; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_181 = _inst_type_T_13 ? 3'h1 : _inst_type_T_180; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_182 = _inst_type_T_11 ? 3'h1 : _inst_type_T_181; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_183 = _inst_type_T_9 ? 3'h1 : _inst_type_T_182; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_184 = _inst_type_T_7 ? 3'h2 : _inst_type_T_183; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_185 = _inst_type_T_5 ? 3'h1 : _inst_type_T_184; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_186 = _inst_type_T_3 ? 3'h3 : _inst_type_T_185; // @[Lookup.scala 33:37]
  wire [2:0] inst_type_2 = _inst_type_T_1 ? 3'h2 : _inst_type_T_186; // @[Lookup.scala 33:37]
  wire  _inst_type_T_235 = _inst_type_T_53 ? 1'h0 : _inst_type_T_55 | (_inst_type_T_57 | (_inst_type_T_59 | (
    _inst_type_T_61 | (_inst_type_T_63 | (_inst_type_T_65 | (_inst_type_T_67 | (_inst_type_T_69 | (_inst_type_T_71 |
    _inst_type_T_73)))))))); // @[Lookup.scala 33:37]
  wire  _inst_type_T_236 = _inst_type_T_51 ? 1'h0 : _inst_type_T_235; // @[Lookup.scala 33:37]
  wire  _inst_type_T_237 = _inst_type_T_49 ? 1'h0 : _inst_type_T_236; // @[Lookup.scala 33:37]
  wire  _inst_type_T_238 = _inst_type_T_47 ? 1'h0 : _inst_type_T_237; // @[Lookup.scala 33:37]
  wire  _inst_type_T_239 = _inst_type_T_45 ? 1'h0 : _inst_type_T_238; // @[Lookup.scala 33:37]
  wire  _inst_type_T_240 = _inst_type_T_43 ? 1'h0 : _inst_type_T_239; // @[Lookup.scala 33:37]
  wire  _inst_type_T_260 = _inst_type_T_3 ? 1'h0 : _inst_type_T_5 | (_inst_type_T_7 | (_inst_type_T_9 | (_inst_type_T_11
     | (_inst_type_T_13 | (_inst_type_T_15 | (_inst_type_T_17 | (_inst_type_T_19 | (_inst_type_T_21 | (_inst_type_T_23
     | (_inst_type_T_25 | (_inst_type_T_27 | (_inst_type_T_29 | (_inst_type_T_31 | (_inst_type_T_33 | (_inst_type_T_35
     | (_inst_type_T_37 | (_inst_type_T_39 | (_inst_type_T_41 | _inst_type_T_240)))))))))))))))))); // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_262 = _inst_type_T_73 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_263 = _inst_type_T_71 ? 3'h3 : _inst_type_T_262; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_264 = _inst_type_T_69 ? 3'h3 : _inst_type_T_263; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_265 = _inst_type_T_67 ? 3'h3 : _inst_type_T_264; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_266 = _inst_type_T_65 ? 3'h3 : _inst_type_T_265; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_267 = _inst_type_T_63 ? 3'h3 : _inst_type_T_266; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_268 = _inst_type_T_61 ? 3'h0 : _inst_type_T_267; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_269 = _inst_type_T_59 ? 3'h0 : _inst_type_T_268; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_270 = _inst_type_T_57 ? 3'h2 : _inst_type_T_269; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_271 = _inst_type_T_55 ? 3'h2 : _inst_type_T_270; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_272 = _inst_type_T_53 ? 3'h0 : _inst_type_T_271; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_273 = _inst_type_T_51 ? 3'h0 : _inst_type_T_272; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_274 = _inst_type_T_49 ? 3'h0 : _inst_type_T_273; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_275 = _inst_type_T_47 ? 3'h0 : _inst_type_T_274; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_276 = _inst_type_T_45 ? 3'h0 : _inst_type_T_275; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_277 = _inst_type_T_43 ? 3'h0 : _inst_type_T_276; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_278 = _inst_type_T_41 ? 3'h0 : _inst_type_T_277; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_279 = _inst_type_T_39 ? 3'h0 : _inst_type_T_278; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_280 = _inst_type_T_37 ? 3'h0 : _inst_type_T_279; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_281 = _inst_type_T_35 ? 3'h0 : _inst_type_T_280; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_282 = _inst_type_T_33 ? 3'h0 : _inst_type_T_281; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_283 = _inst_type_T_31 ? 3'h0 : _inst_type_T_282; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_284 = _inst_type_T_29 ? 3'h0 : _inst_type_T_283; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_285 = _inst_type_T_27 ? 3'h0 : _inst_type_T_284; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_286 = _inst_type_T_25 ? 3'h0 : _inst_type_T_285; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_287 = _inst_type_T_23 ? 3'h0 : _inst_type_T_286; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_288 = _inst_type_T_21 ? 3'h0 : _inst_type_T_287; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_289 = _inst_type_T_19 ? 3'h0 : _inst_type_T_288; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_290 = _inst_type_T_17 ? 3'h0 : _inst_type_T_289; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_291 = _inst_type_T_15 ? 3'h0 : _inst_type_T_290; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_292 = _inst_type_T_13 ? 3'h0 : _inst_type_T_291; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_293 = _inst_type_T_11 ? 3'h0 : _inst_type_T_292; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_294 = _inst_type_T_9 ? 3'h0 : _inst_type_T_293; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_295 = _inst_type_T_7 ? 3'h0 : _inst_type_T_294; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_296 = _inst_type_T_5 ? 3'h0 : _inst_type_T_295; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_297 = _inst_type_T_3 ? 3'h0 : _inst_type_T_296; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_298 = _inst_type_T_75 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_299 = _inst_type_T_73 ? 3'h3 : _inst_type_T_298; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_300 = _inst_type_T_71 ? 3'h3 : _inst_type_T_299; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_301 = _inst_type_T_69 ? 3'h2 : _inst_type_T_300; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_302 = _inst_type_T_67 ? 3'h2 : _inst_type_T_301; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_303 = _inst_type_T_65 ? 3'h1 : _inst_type_T_302; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_304 = _inst_type_T_63 ? 3'h1 : _inst_type_T_303; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_305 = _inst_type_T_61 ? 3'h0 : _inst_type_T_304; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_306 = _inst_type_T_59 ? 3'h0 : _inst_type_T_305; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_307 = _inst_type_T_57 ? 3'h0 : _inst_type_T_306; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_308 = _inst_type_T_55 ? 3'h0 : _inst_type_T_307; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_309 = _inst_type_T_53 ? 3'h0 : _inst_type_T_308; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_310 = _inst_type_T_51 ? 3'h0 : _inst_type_T_309; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_311 = _inst_type_T_49 ? 3'h0 : _inst_type_T_310; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_312 = _inst_type_T_47 ? 3'h0 : _inst_type_T_311; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_313 = _inst_type_T_45 ? 3'h0 : _inst_type_T_312; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_314 = _inst_type_T_43 ? 3'h0 : _inst_type_T_313; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_315 = _inst_type_T_41 ? 3'h0 : _inst_type_T_314; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_316 = _inst_type_T_39 ? 3'h0 : _inst_type_T_315; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_317 = _inst_type_T_37 ? 3'h0 : _inst_type_T_316; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_318 = _inst_type_T_35 ? 3'h0 : _inst_type_T_317; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_319 = _inst_type_T_33 ? 3'h0 : _inst_type_T_318; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_320 = _inst_type_T_31 ? 3'h0 : _inst_type_T_319; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_321 = _inst_type_T_29 ? 3'h0 : _inst_type_T_320; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_322 = _inst_type_T_27 ? 3'h0 : _inst_type_T_321; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_323 = _inst_type_T_25 ? 3'h0 : _inst_type_T_322; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_324 = _inst_type_T_23 ? 3'h0 : _inst_type_T_323; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_325 = _inst_type_T_21 ? 3'h0 : _inst_type_T_324; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_326 = _inst_type_T_19 ? 3'h0 : _inst_type_T_325; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_327 = _inst_type_T_17 ? 3'h0 : _inst_type_T_326; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_328 = _inst_type_T_15 ? 3'h0 : _inst_type_T_327; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_329 = _inst_type_T_13 ? 3'h0 : _inst_type_T_328; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_330 = _inst_type_T_11 ? 3'h0 : _inst_type_T_329; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_331 = _inst_type_T_9 ? 3'h0 : _inst_type_T_330; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_332 = _inst_type_T_7 ? 3'h0 : _inst_type_T_331; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_333 = _inst_type_T_5 ? 3'h0 : _inst_type_T_332; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_334 = _inst_type_T_3 ? 3'h0 : _inst_type_T_333; // @[Lookup.scala 33:37]
  wire  _op1_data_T = inst_type_1 == 2'h0; // @[ID.scala 168:18]
  wire  _op1_data_T_1 = inst_type_1 == 2'h1; // @[ID.scala 169:18]
  wire  _op1_data_T_2 = inst_type_1 == 2'h3; // @[ID.scala 170:18]
  wire [31:0] _op1_data_T_3 = _op1_data_T_2 ? imm_z_uext : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _op1_data_T_4 = _op1_data_T_1 ? io_in_if_in_reg_pc : _op1_data_T_3; // @[Mux.scala 98:16]
  wire [31:0] op1_data = _op1_data_T ? rs1_data : _op1_data_T_4; // @[Mux.scala 98:16]
  wire  _op2_data_T = inst_type_2 == 3'h1; // @[ID.scala 174:18]
  wire  _op2_data_T_1 = inst_type_2 == 3'h2; // @[ID.scala 175:18]
  wire  _op2_data_T_2 = inst_type_2 == 3'h3; // @[ID.scala 176:18]
  wire  _op2_data_T_3 = inst_type_2 == 3'h4; // @[ID.scala 177:18]
  wire  _op2_data_T_4 = inst_type_2 == 3'h5; // @[ID.scala 178:18]
  wire [31:0] _op2_data_T_5 = _op2_data_T_4 ? imm_u_shifted : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_6 = _op2_data_T_3 ? imm_j_sext : _op2_data_T_5; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_7 = _op2_data_T_2 ? imm_s_sext : _op2_data_T_6; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_8 = _op2_data_T_1 ? imm_i_sext : _op2_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] op2_data = _op2_data_T ? rs2_data : _op2_data_T_8; // @[Mux.scala 98:16]
  wire [31:0] _GEN_128 = {{27'd0}, io_in_wb_in_rd_addr}; // @[ID.scala 182:45]
  wire  _T_4 = ~reset; // @[ID.scala 202:11]
  assign io_out_op1_data = _op1_data_T ? rs1_data : _op1_data_T_4; // @[Mux.scala 98:16]
  assign io_out_op2_data = _op2_data_T ? rs2_data : _op2_data_T_8; // @[Mux.scala 98:16]
  assign io_out_rd_addr = inst[11:7]; // @[ID.scala 97:24]
  assign io_out_csr_addr_default = {{20'd0}, csr_addr_default}; // @[ID.scala 98:32]
  assign io_out_exe_fun = _inst_type_T_1 ? 5'h1 : _inst_type_T_112; // @[Lookup.scala 33:37]
  assign io_out_mem_wen = _inst_type_T_1 ? 1'h0 : _inst_type_T_3; // @[Lookup.scala 33:37]
  assign io_out_rd_wen = _inst_type_T_1 | _inst_type_T_260; // @[Lookup.scala 33:37]
  assign io_out_rd_sel = _inst_type_T_1 ? 3'h1 : _inst_type_T_297; // @[Lookup.scala 33:37]
  assign io_out_csr_cmd = _inst_type_T_1 ? 3'h0 : _inst_type_T_334; // @[Lookup.scala 33:37]
  assign io_out_rs2_data = _rs2_data_T ? 32'h0 : _rs2_data_T_8; // @[Mux.scala 98:16]
  assign io_out_imm_b_sext = {imm_b_sext_hi,1'h0}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[ID.scala 75:26]
      reg_x_0 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h0 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_0 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_1 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_1 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_2 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h2 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_2 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_3 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h3 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_3 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_4 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h4 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_4 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_5 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h5 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_5 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_6 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h6 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_6 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_7 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h7 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_7 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_8 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h8 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_8 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_9 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h9 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_9 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_10 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'ha == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_10 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_11 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hb == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_11 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_12 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hc == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_12 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_13 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hd == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_13 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_14 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'he == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_14 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_15 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hf == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_15 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_16 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h10 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_16 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_17 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h11 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_17 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_18 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h12 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_18 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_19 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h13 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_19 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_20 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h14 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_20 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_21 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h15 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_21 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_22 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h16 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_22 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_23 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h17 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_23 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_24 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h18 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_24 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_25 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h19 == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_25 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_26 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1a == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_26 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_27 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1b == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_27 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_28 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1c == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_28 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_29 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1d == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_29 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_30 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1e == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_30 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_31 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_in_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1f == io_in_wb_in_rd_addr) begin // @[ID.scala 183:27]
        reg_x_31 <= io_in_wb_in_rd_data; // @[ID.scala 183:27]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------ID------------\n"); // @[ID.scala 202:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"rs1_addr: %d\n",rs1_addr); // @[ID.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"rs2_addr: %d\n",rs2_addr); // @[ID.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"op1_data: 0x%x\n",op1_data); // @[ID.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"op2_data: 0x%x\n",op2_data); // @[ID.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"stall_flag: %d\n",io_in_stall_in_stall_flag); // @[ID.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_x_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_x_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_x_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_x_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_x_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_x_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_x_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_x_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_x_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_x_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_x_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_x_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_x_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_x_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_x_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_x_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_x_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_x_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_x_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_x_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_x_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_x_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_x_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_x_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_x_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_x_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_x_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_x_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_x_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_x_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_x_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_x_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stall(
  input  [31:0] io_in_if_in_inst,
  input  [4:0]  io_in_id_reg_in_rd_addr,
  input         io_in_id_reg_in_rd_wen,
  output        io_out_stall_flag
);
  wire [4:0] rs1_addr_default = io_in_if_in_inst[19:15]; // @[Stall.scala 27:43]
  wire [4:0] rs2_addr_default = io_in_if_in_inst[24:20]; // @[Stall.scala 28:43]
  wire  rs1_data_hazard = io_in_id_reg_in_rd_wen & rs1_addr_default != 5'h0 & rs1_addr_default ==
    io_in_id_reg_in_rd_addr; // @[Stall.scala 29:84]
  wire  rs2_data_hazard = io_in_id_reg_in_rd_wen & rs2_addr_default != 5'h0 & rs2_addr_default ==
    io_in_id_reg_in_rd_addr; // @[Stall.scala 30:84]
  assign io_out_stall_flag = rs1_data_hazard | rs2_data_hazard; // @[Stall.scala 31:39]
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_in_id_in_op1_data,
  input  [31:0] io_in_id_in_op2_data,
  input  [4:0]  io_in_id_in_exe_fun,
  input  [2:0]  io_in_id_in_rd_sel,
  output [31:0] io_out_alu_out,
  output        io_out_jump_flag
);
  wire  _alu_out_T = io_in_id_in_exe_fun == 5'h1; // @[ALU.scala 55:18]
  wire [31:0] _alu_out_T_2 = io_in_id_in_op1_data + io_in_id_in_op2_data; // @[ALU.scala 55:46]
  wire  _alu_out_T_3 = io_in_id_in_exe_fun == 5'h2; // @[ALU.scala 56:18]
  wire [31:0] _alu_out_T_5 = io_in_id_in_op1_data - io_in_id_in_op2_data; // @[ALU.scala 56:46]
  wire  _alu_out_T_6 = io_in_id_in_exe_fun == 5'h3; // @[ALU.scala 57:18]
  wire [31:0] _alu_out_T_7 = io_in_id_in_op1_data & io_in_id_in_op2_data; // @[ALU.scala 57:46]
  wire  _alu_out_T_8 = io_in_id_in_exe_fun == 5'h4; // @[ALU.scala 58:18]
  wire [31:0] _alu_out_T_9 = io_in_id_in_op1_data | io_in_id_in_op2_data; // @[ALU.scala 58:46]
  wire  _alu_out_T_10 = io_in_id_in_exe_fun == 5'h5; // @[ALU.scala 59:18]
  wire [31:0] _alu_out_T_11 = io_in_id_in_op1_data ^ io_in_id_in_op2_data; // @[ALU.scala 59:46]
  wire  _alu_out_T_12 = io_in_id_in_exe_fun == 5'h6; // @[ALU.scala 60:18]
  wire [62:0] _GEN_0 = {{31'd0}, io_in_id_in_op1_data}; // @[ALU.scala 60:46]
  wire [62:0] _alu_out_T_14 = _GEN_0 << io_in_id_in_op2_data[4:0]; // @[ALU.scala 60:46]
  wire  _alu_out_T_16 = io_in_id_in_exe_fun == 5'h7; // @[ALU.scala 61:18]
  wire [31:0] _alu_out_T_18 = io_in_id_in_op1_data >> io_in_id_in_op2_data[4:0]; // @[ALU.scala 61:46]
  wire  _alu_out_T_19 = io_in_id_in_exe_fun == 5'h8; // @[ALU.scala 62:18]
  wire [31:0] _alu_out_T_23 = $signed(io_in_id_in_op1_data) >>> io_in_id_in_op2_data[4:0]; // @[ALU.scala 62:80]
  wire  _alu_out_T_24 = io_in_id_in_exe_fun == 5'h9; // @[ALU.scala 63:18]
  wire  _alu_out_T_27 = $signed(io_in_id_in_op1_data) < $signed(io_in_id_in_op2_data); // @[ALU.scala 63:55]
  wire  _alu_out_T_28 = io_in_id_in_exe_fun == 5'ha; // @[ALU.scala 64:18]
  wire  _alu_out_T_29 = io_in_id_in_op1_data < io_in_id_in_op2_data; // @[ALU.scala 64:46]
  wire  _alu_out_T_30 = io_in_id_in_exe_fun == 5'h11; // @[ALU.scala 65:18]
  wire [31:0] _alu_out_T_34 = _alu_out_T_2 & 32'hfffffffe; // @[ALU.scala 65:59]
  wire  _alu_out_T_35 = io_in_id_in_exe_fun == 5'h12; // @[ALU.scala 66:18]
  wire [31:0] _alu_out_T_36 = _alu_out_T_35 ? io_in_id_in_op1_data : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_37 = _alu_out_T_30 ? _alu_out_T_34 : _alu_out_T_36; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_38 = _alu_out_T_28 ? {{31'd0}, _alu_out_T_29} : _alu_out_T_37; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_39 = _alu_out_T_24 ? {{31'd0}, _alu_out_T_27} : _alu_out_T_38; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_40 = _alu_out_T_19 ? _alu_out_T_23 : _alu_out_T_39; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_41 = _alu_out_T_16 ? _alu_out_T_18 : _alu_out_T_40; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_42 = _alu_out_T_12 ? _alu_out_T_14[31:0] : _alu_out_T_41; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_43 = _alu_out_T_10 ? _alu_out_T_11 : _alu_out_T_42; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_44 = _alu_out_T_8 ? _alu_out_T_9 : _alu_out_T_43; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_45 = _alu_out_T_6 ? _alu_out_T_7 : _alu_out_T_44; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_46 = _alu_out_T_3 ? _alu_out_T_5 : _alu_out_T_45; // @[Mux.scala 98:16]
  wire [31:0] alu_out = _alu_out_T ? _alu_out_T_2 : _alu_out_T_46; // @[Mux.scala 98:16]
  wire  jump_flag = io_in_id_in_rd_sel == 3'h2; // @[ALU.scala 69:29]
  wire  _T_1 = ~reset; // @[ALU.scala 76:11]
  assign io_out_alu_out = _alu_out_T ? _alu_out_T_2 : _alu_out_T_46; // @[Mux.scala 98:16]
  assign io_out_jump_flag = io_in_id_in_rd_sel == 3'h2; // @[ALU.scala 69:29]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------EX------------\n"); // @[ALU.scala 76:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"alu_out: 0x%x\n",alu_out); // @[ALU.scala 77:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"jump_flg: %d\n",jump_flag); // @[ALU.scala 78:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BR(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_in_reg_pc,
  input  [31:0] io_in_id_in_op1_data,
  input  [31:0] io_in_id_in_op2_data,
  input  [4:0]  io_in_id_in_exe_fun,
  input  [31:0] io_in_id_in_imm_b_sext,
  output        io_out_br_flag,
  output [31:0] io_out_br_target
);
  wire [31:0] br_target = io_in_if_in_reg_pc + io_in_id_in_imm_b_sext; // @[BR.scala 56:30]
  wire  _br_flag_T = io_in_id_in_exe_fun == 5'hb; // @[BR.scala 58:18]
  wire  _br_flag_T_1 = io_in_id_in_op1_data == io_in_id_in_op2_data; // @[BR.scala 58:45]
  wire  _br_flag_T_2 = io_in_id_in_exe_fun == 5'hc; // @[BR.scala 59:18]
  wire  _br_flag_T_4 = ~_br_flag_T_1; // @[BR.scala 59:34]
  wire  _br_flag_T_5 = io_in_id_in_exe_fun == 5'hd; // @[BR.scala 60:18]
  wire  _br_flag_T_8 = $signed(io_in_id_in_op1_data) < $signed(io_in_id_in_op2_data); // @[BR.scala 60:54]
  wire  _br_flag_T_9 = io_in_id_in_exe_fun == 5'he; // @[BR.scala 61:18]
  wire  _br_flag_T_13 = ~_br_flag_T_8; // @[BR.scala 61:34]
  wire  _br_flag_T_14 = io_in_id_in_exe_fun == 5'hf; // @[BR.scala 62:18]
  wire  _br_flag_T_15 = io_in_id_in_op1_data < io_in_id_in_op2_data; // @[BR.scala 62:45]
  wire  _br_flag_T_16 = io_in_id_in_exe_fun == 5'h10; // @[BR.scala 63:18]
  wire  _br_flag_T_18 = ~_br_flag_T_15; // @[BR.scala 63:34]
  wire  _br_flag_T_20 = _br_flag_T_14 ? _br_flag_T_15 : _br_flag_T_16 & _br_flag_T_18; // @[Mux.scala 98:16]
  wire  _br_flag_T_21 = _br_flag_T_9 ? _br_flag_T_13 : _br_flag_T_20; // @[Mux.scala 98:16]
  wire  _br_flag_T_22 = _br_flag_T_5 ? _br_flag_T_8 : _br_flag_T_21; // @[Mux.scala 98:16]
  wire  _br_flag_T_23 = _br_flag_T_2 ? _br_flag_T_4 : _br_flag_T_22; // @[Mux.scala 98:16]
  wire  br_flag = _br_flag_T ? _br_flag_T_1 : _br_flag_T_23; // @[Mux.scala 98:16]
  wire  _T_1 = ~reset; // @[BR.scala 71:11]
  assign io_out_br_flag = _br_flag_T ? _br_flag_T_1 : _br_flag_T_23; // @[Mux.scala 98:16]
  assign io_out_br_target = io_in_if_in_reg_pc + io_in_id_in_imm_b_sext; // @[BR.scala 56:30]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"branch_flg: %d\n",br_flag); // @[BR.scala 71:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"branch_target: 0x%x\n",br_target); // @[BR.scala 72:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MEM(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_in_reg_pc,
  input  [31:0] io_in_id_in_op1_data,
  input  [4:0]  io_in_id_in_rd_addr,
  input  [31:0] io_in_id_in_csr_addr_default,
  input         io_in_id_in_mem_wen,
  input         io_in_id_in_rd_wen,
  input  [2:0]  io_in_id_in_rd_sel,
  input  [2:0]  io_in_id_in_csr_cmd,
  input  [31:0] io_in_id_in_rs2_data,
  input  [31:0] io_in_ex_in_alu_out,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data,
  output [31:0] io_datamem_addr,
  input  [31:0] io_datamem_rdata,
  output        io_datamem_wen,
  output [31:0] io_datamem_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_csr_0; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_2; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_3; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_4; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_5; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_6; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_7; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_8; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_9; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_10; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_11; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_12; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_13; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_14; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_15; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_16; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_17; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_18; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_19; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_20; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_21; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_22; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_23; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_24; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_25; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_26; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_27; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_28; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_29; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_30; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_31; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_32; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_33; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_34; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_35; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_36; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_37; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_38; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_39; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_40; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_41; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_42; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_43; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_44; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_45; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_46; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_47; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_48; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_49; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_50; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_51; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_52; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_53; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_54; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_55; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_56; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_57; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_58; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_59; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_60; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_61; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_62; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_63; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_64; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_65; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_66; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_67; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_68; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_69; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_70; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_71; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_72; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_73; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_74; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_75; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_76; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_77; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_78; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_79; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_80; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_81; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_82; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_83; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_84; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_85; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_86; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_87; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_88; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_89; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_90; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_91; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_92; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_93; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_94; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_95; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_96; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_97; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_98; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_99; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_100; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_101; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_102; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_103; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_104; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_105; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_106; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_107; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_108; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_109; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_110; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_111; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_112; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_113; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_114; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_115; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_116; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_117; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_118; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_119; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_120; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_121; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_122; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_123; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_124; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_125; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_126; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_127; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_128; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_129; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_130; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_131; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_132; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_133; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_134; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_135; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_136; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_137; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_138; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_139; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_140; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_141; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_142; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_143; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_144; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_145; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_146; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_147; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_148; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_149; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_150; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_151; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_152; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_153; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_154; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_155; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_156; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_157; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_158; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_159; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_160; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_161; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_162; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_163; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_164; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_165; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_166; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_167; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_168; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_169; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_170; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_171; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_172; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_173; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_174; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_175; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_176; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_177; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_178; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_179; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_180; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_181; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_182; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_183; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_184; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_185; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_186; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_187; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_188; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_189; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_190; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_191; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_192; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_193; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_194; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_195; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_196; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_197; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_198; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_199; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_200; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_201; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_202; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_203; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_204; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_205; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_206; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_207; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_208; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_209; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_210; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_211; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_212; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_213; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_214; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_215; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_216; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_217; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_218; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_219; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_220; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_221; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_222; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_223; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_224; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_225; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_226; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_227; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_228; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_229; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_230; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_231; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_232; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_233; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_234; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_235; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_236; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_237; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_238; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_239; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_240; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_241; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_242; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_243; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_244; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_245; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_246; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_247; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_248; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_249; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_250; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_251; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_252; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_253; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_254; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_255; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_256; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_257; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_258; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_259; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_260; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_261; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_262; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_263; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_264; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_265; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_266; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_267; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_268; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_269; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_270; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_271; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_272; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_273; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_274; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_275; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_276; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_277; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_278; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_279; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_280; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_281; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_282; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_283; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_284; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_285; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_286; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_287; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_288; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_289; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_290; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_291; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_292; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_293; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_294; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_295; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_296; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_297; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_298; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_299; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_300; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_301; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_302; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_303; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_304; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_305; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_306; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_307; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_308; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_309; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_310; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_311; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_312; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_313; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_314; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_315; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_316; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_317; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_318; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_319; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_320; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_321; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_322; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_323; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_324; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_325; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_326; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_327; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_328; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_329; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_330; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_331; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_332; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_333; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_334; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_335; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_336; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_337; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_338; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_339; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_340; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_341; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_342; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_343; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_344; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_345; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_346; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_347; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_348; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_349; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_350; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_351; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_352; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_353; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_354; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_355; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_356; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_357; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_358; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_359; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_360; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_361; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_362; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_363; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_364; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_365; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_366; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_367; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_368; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_369; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_370; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_371; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_372; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_373; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_374; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_375; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_376; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_377; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_378; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_379; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_380; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_381; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_382; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_383; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_384; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_385; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_386; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_387; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_388; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_389; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_390; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_391; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_392; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_393; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_394; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_395; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_396; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_397; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_398; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_399; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_400; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_401; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_402; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_403; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_404; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_405; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_406; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_407; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_408; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_409; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_410; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_411; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_412; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_413; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_414; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_415; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_416; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_417; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_418; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_419; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_420; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_421; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_422; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_423; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_424; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_425; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_426; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_427; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_428; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_429; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_430; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_431; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_432; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_433; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_434; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_435; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_436; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_437; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_438; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_439; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_440; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_441; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_442; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_443; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_444; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_445; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_446; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_447; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_448; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_449; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_450; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_451; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_452; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_453; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_454; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_455; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_456; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_457; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_458; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_459; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_460; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_461; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_462; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_463; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_464; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_465; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_466; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_467; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_468; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_469; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_470; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_471; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_472; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_473; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_474; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_475; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_476; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_477; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_478; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_479; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_480; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_481; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_482; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_483; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_484; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_485; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_486; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_487; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_488; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_489; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_490; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_491; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_492; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_493; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_494; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_495; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_496; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_497; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_498; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_499; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_500; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_501; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_502; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_503; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_504; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_505; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_506; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_507; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_508; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_509; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_510; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_511; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_512; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_513; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_514; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_515; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_516; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_517; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_518; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_519; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_520; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_521; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_522; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_523; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_524; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_525; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_526; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_527; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_528; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_529; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_530; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_531; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_532; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_533; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_534; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_535; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_536; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_537; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_538; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_539; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_540; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_541; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_542; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_543; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_544; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_545; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_546; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_547; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_548; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_549; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_550; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_551; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_552; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_553; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_554; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_555; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_556; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_557; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_558; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_559; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_560; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_561; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_562; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_563; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_564; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_565; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_566; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_567; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_568; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_569; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_570; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_571; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_572; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_573; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_574; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_575; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_576; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_577; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_578; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_579; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_580; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_581; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_582; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_583; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_584; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_585; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_586; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_587; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_588; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_589; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_590; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_591; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_592; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_593; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_594; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_595; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_596; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_597; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_598; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_599; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_600; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_601; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_602; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_603; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_604; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_605; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_606; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_607; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_608; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_609; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_610; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_611; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_612; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_613; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_614; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_615; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_616; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_617; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_618; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_619; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_620; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_621; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_622; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_623; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_624; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_625; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_626; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_627; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_628; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_629; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_630; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_631; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_632; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_633; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_634; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_635; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_636; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_637; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_638; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_639; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_640; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_641; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_642; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_643; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_644; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_645; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_646; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_647; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_648; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_649; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_650; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_651; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_652; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_653; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_654; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_655; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_656; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_657; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_658; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_659; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_660; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_661; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_662; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_663; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_664; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_665; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_666; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_667; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_668; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_669; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_670; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_671; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_672; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_673; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_674; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_675; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_676; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_677; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_678; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_679; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_680; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_681; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_682; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_683; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_684; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_685; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_686; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_687; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_688; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_689; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_690; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_691; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_692; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_693; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_694; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_695; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_696; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_697; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_698; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_699; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_700; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_701; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_702; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_703; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_704; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_705; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_706; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_707; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_708; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_709; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_710; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_711; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_712; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_713; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_714; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_715; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_716; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_717; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_718; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_719; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_720; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_721; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_722; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_723; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_724; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_725; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_726; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_727; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_728; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_729; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_730; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_731; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_732; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_733; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_734; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_735; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_736; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_737; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_738; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_739; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_740; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_741; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_742; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_743; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_744; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_745; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_746; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_747; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_748; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_749; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_750; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_751; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_752; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_753; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_754; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_755; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_756; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_757; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_758; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_759; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_760; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_761; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_762; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_763; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_764; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_765; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_766; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_767; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_768; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_769; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_770; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_771; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_772; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_773; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_774; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_775; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_776; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_777; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_778; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_779; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_780; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_781; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_782; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_783; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_784; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_785; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_786; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_787; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_788; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_789; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_790; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_791; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_792; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_793; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_794; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_795; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_796; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_797; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_798; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_799; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_800; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_801; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_802; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_803; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_804; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_805; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_806; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_807; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_808; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_809; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_810; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_811; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_812; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_813; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_814; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_815; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_816; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_817; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_818; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_819; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_820; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_821; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_822; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_823; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_824; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_825; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_826; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_827; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_828; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_829; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_830; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_831; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_832; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_833; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_834; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_835; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_836; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_837; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_838; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_839; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_840; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_841; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_842; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_843; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_844; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_845; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_846; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_847; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_848; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_849; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_850; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_851; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_852; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_853; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_854; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_855; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_856; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_857; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_858; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_859; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_860; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_861; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_862; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_863; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_864; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_865; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_866; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_867; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_868; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_869; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_870; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_871; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_872; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_873; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_874; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_875; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_876; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_877; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_878; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_879; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_880; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_881; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_882; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_883; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_884; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_885; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_886; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_887; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_888; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_889; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_890; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_891; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_892; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_893; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_894; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_895; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_896; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_897; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_898; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_899; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_900; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_901; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_902; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_903; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_904; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_905; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_906; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_907; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_908; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_909; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_910; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_911; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_912; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_913; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_914; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_915; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_916; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_917; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_918; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_919; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_920; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_921; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_922; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_923; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_924; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_925; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_926; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_927; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_928; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_929; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_930; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_931; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_932; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_933; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_934; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_935; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_936; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_937; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_938; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_939; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_940; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_941; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_942; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_943; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_944; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_945; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_946; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_947; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_948; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_949; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_950; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_951; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_952; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_953; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_954; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_955; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_956; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_957; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_958; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_959; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_960; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_961; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_962; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_963; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_964; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_965; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_966; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_967; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_968; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_969; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_970; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_971; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_972; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_973; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_974; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_975; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_976; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_977; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_978; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_979; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_980; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_981; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_982; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_983; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_984; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_985; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_986; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_987; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_988; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_989; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_990; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_991; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_992; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_993; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_994; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_995; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_996; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_997; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_998; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_999; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1000; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1001; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1002; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1003; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1004; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1005; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1006; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1007; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1008; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1009; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1010; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1011; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1012; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1013; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1014; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1015; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1016; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1017; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1018; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1019; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1020; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1021; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1022; // @[MEM.scala 54:26]
  reg [31:0] reg_csr_1023; // @[MEM.scala 54:26]
  wire  _csr_addr_T = io_in_id_in_csr_cmd == 3'h4; // @[MEM.scala 78:18]
  wire [31:0] csr_addr = _csr_addr_T ? 32'h342 : io_in_id_in_csr_addr_default; // @[Mux.scala 98:16]
  wire  _csr_wdata_T = io_in_id_in_csr_cmd == 3'h1; // @[MEM.scala 82:18]
  wire  _csr_wdata_T_1 = io_in_id_in_csr_cmd == 3'h2; // @[MEM.scala 83:18]
  wire [31:0] _GEN_1 = 10'h1 == csr_addr[9:0] ? reg_csr_1 : reg_csr_0; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_2 = 10'h2 == csr_addr[9:0] ? reg_csr_2 : _GEN_1; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_3 = 10'h3 == csr_addr[9:0] ? reg_csr_3 : _GEN_2; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_4 = 10'h4 == csr_addr[9:0] ? reg_csr_4 : _GEN_3; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_5 = 10'h5 == csr_addr[9:0] ? reg_csr_5 : _GEN_4; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_6 = 10'h6 == csr_addr[9:0] ? reg_csr_6 : _GEN_5; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_7 = 10'h7 == csr_addr[9:0] ? reg_csr_7 : _GEN_6; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_8 = 10'h8 == csr_addr[9:0] ? reg_csr_8 : _GEN_7; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_9 = 10'h9 == csr_addr[9:0] ? reg_csr_9 : _GEN_8; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_10 = 10'ha == csr_addr[9:0] ? reg_csr_10 : _GEN_9; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_11 = 10'hb == csr_addr[9:0] ? reg_csr_11 : _GEN_10; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_12 = 10'hc == csr_addr[9:0] ? reg_csr_12 : _GEN_11; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_13 = 10'hd == csr_addr[9:0] ? reg_csr_13 : _GEN_12; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_14 = 10'he == csr_addr[9:0] ? reg_csr_14 : _GEN_13; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_15 = 10'hf == csr_addr[9:0] ? reg_csr_15 : _GEN_14; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_16 = 10'h10 == csr_addr[9:0] ? reg_csr_16 : _GEN_15; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_17 = 10'h11 == csr_addr[9:0] ? reg_csr_17 : _GEN_16; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_18 = 10'h12 == csr_addr[9:0] ? reg_csr_18 : _GEN_17; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_19 = 10'h13 == csr_addr[9:0] ? reg_csr_19 : _GEN_18; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_20 = 10'h14 == csr_addr[9:0] ? reg_csr_20 : _GEN_19; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_21 = 10'h15 == csr_addr[9:0] ? reg_csr_21 : _GEN_20; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_22 = 10'h16 == csr_addr[9:0] ? reg_csr_22 : _GEN_21; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_23 = 10'h17 == csr_addr[9:0] ? reg_csr_23 : _GEN_22; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_24 = 10'h18 == csr_addr[9:0] ? reg_csr_24 : _GEN_23; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_25 = 10'h19 == csr_addr[9:0] ? reg_csr_25 : _GEN_24; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_26 = 10'h1a == csr_addr[9:0] ? reg_csr_26 : _GEN_25; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_27 = 10'h1b == csr_addr[9:0] ? reg_csr_27 : _GEN_26; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_28 = 10'h1c == csr_addr[9:0] ? reg_csr_28 : _GEN_27; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_29 = 10'h1d == csr_addr[9:0] ? reg_csr_29 : _GEN_28; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_30 = 10'h1e == csr_addr[9:0] ? reg_csr_30 : _GEN_29; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_31 = 10'h1f == csr_addr[9:0] ? reg_csr_31 : _GEN_30; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_32 = 10'h20 == csr_addr[9:0] ? reg_csr_32 : _GEN_31; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_33 = 10'h21 == csr_addr[9:0] ? reg_csr_33 : _GEN_32; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_34 = 10'h22 == csr_addr[9:0] ? reg_csr_34 : _GEN_33; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_35 = 10'h23 == csr_addr[9:0] ? reg_csr_35 : _GEN_34; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_36 = 10'h24 == csr_addr[9:0] ? reg_csr_36 : _GEN_35; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_37 = 10'h25 == csr_addr[9:0] ? reg_csr_37 : _GEN_36; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_38 = 10'h26 == csr_addr[9:0] ? reg_csr_38 : _GEN_37; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_39 = 10'h27 == csr_addr[9:0] ? reg_csr_39 : _GEN_38; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_40 = 10'h28 == csr_addr[9:0] ? reg_csr_40 : _GEN_39; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_41 = 10'h29 == csr_addr[9:0] ? reg_csr_41 : _GEN_40; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_42 = 10'h2a == csr_addr[9:0] ? reg_csr_42 : _GEN_41; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_43 = 10'h2b == csr_addr[9:0] ? reg_csr_43 : _GEN_42; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_44 = 10'h2c == csr_addr[9:0] ? reg_csr_44 : _GEN_43; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_45 = 10'h2d == csr_addr[9:0] ? reg_csr_45 : _GEN_44; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_46 = 10'h2e == csr_addr[9:0] ? reg_csr_46 : _GEN_45; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_47 = 10'h2f == csr_addr[9:0] ? reg_csr_47 : _GEN_46; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_48 = 10'h30 == csr_addr[9:0] ? reg_csr_48 : _GEN_47; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_49 = 10'h31 == csr_addr[9:0] ? reg_csr_49 : _GEN_48; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_50 = 10'h32 == csr_addr[9:0] ? reg_csr_50 : _GEN_49; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_51 = 10'h33 == csr_addr[9:0] ? reg_csr_51 : _GEN_50; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_52 = 10'h34 == csr_addr[9:0] ? reg_csr_52 : _GEN_51; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_53 = 10'h35 == csr_addr[9:0] ? reg_csr_53 : _GEN_52; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_54 = 10'h36 == csr_addr[9:0] ? reg_csr_54 : _GEN_53; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_55 = 10'h37 == csr_addr[9:0] ? reg_csr_55 : _GEN_54; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_56 = 10'h38 == csr_addr[9:0] ? reg_csr_56 : _GEN_55; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_57 = 10'h39 == csr_addr[9:0] ? reg_csr_57 : _GEN_56; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_58 = 10'h3a == csr_addr[9:0] ? reg_csr_58 : _GEN_57; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_59 = 10'h3b == csr_addr[9:0] ? reg_csr_59 : _GEN_58; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_60 = 10'h3c == csr_addr[9:0] ? reg_csr_60 : _GEN_59; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_61 = 10'h3d == csr_addr[9:0] ? reg_csr_61 : _GEN_60; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_62 = 10'h3e == csr_addr[9:0] ? reg_csr_62 : _GEN_61; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_63 = 10'h3f == csr_addr[9:0] ? reg_csr_63 : _GEN_62; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_64 = 10'h40 == csr_addr[9:0] ? reg_csr_64 : _GEN_63; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_65 = 10'h41 == csr_addr[9:0] ? reg_csr_65 : _GEN_64; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_66 = 10'h42 == csr_addr[9:0] ? reg_csr_66 : _GEN_65; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_67 = 10'h43 == csr_addr[9:0] ? reg_csr_67 : _GEN_66; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_68 = 10'h44 == csr_addr[9:0] ? reg_csr_68 : _GEN_67; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_69 = 10'h45 == csr_addr[9:0] ? reg_csr_69 : _GEN_68; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_70 = 10'h46 == csr_addr[9:0] ? reg_csr_70 : _GEN_69; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_71 = 10'h47 == csr_addr[9:0] ? reg_csr_71 : _GEN_70; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_72 = 10'h48 == csr_addr[9:0] ? reg_csr_72 : _GEN_71; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_73 = 10'h49 == csr_addr[9:0] ? reg_csr_73 : _GEN_72; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_74 = 10'h4a == csr_addr[9:0] ? reg_csr_74 : _GEN_73; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_75 = 10'h4b == csr_addr[9:0] ? reg_csr_75 : _GEN_74; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_76 = 10'h4c == csr_addr[9:0] ? reg_csr_76 : _GEN_75; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_77 = 10'h4d == csr_addr[9:0] ? reg_csr_77 : _GEN_76; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_78 = 10'h4e == csr_addr[9:0] ? reg_csr_78 : _GEN_77; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_79 = 10'h4f == csr_addr[9:0] ? reg_csr_79 : _GEN_78; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_80 = 10'h50 == csr_addr[9:0] ? reg_csr_80 : _GEN_79; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_81 = 10'h51 == csr_addr[9:0] ? reg_csr_81 : _GEN_80; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_82 = 10'h52 == csr_addr[9:0] ? reg_csr_82 : _GEN_81; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_83 = 10'h53 == csr_addr[9:0] ? reg_csr_83 : _GEN_82; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_84 = 10'h54 == csr_addr[9:0] ? reg_csr_84 : _GEN_83; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_85 = 10'h55 == csr_addr[9:0] ? reg_csr_85 : _GEN_84; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_86 = 10'h56 == csr_addr[9:0] ? reg_csr_86 : _GEN_85; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_87 = 10'h57 == csr_addr[9:0] ? reg_csr_87 : _GEN_86; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_88 = 10'h58 == csr_addr[9:0] ? reg_csr_88 : _GEN_87; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_89 = 10'h59 == csr_addr[9:0] ? reg_csr_89 : _GEN_88; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_90 = 10'h5a == csr_addr[9:0] ? reg_csr_90 : _GEN_89; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_91 = 10'h5b == csr_addr[9:0] ? reg_csr_91 : _GEN_90; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_92 = 10'h5c == csr_addr[9:0] ? reg_csr_92 : _GEN_91; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_93 = 10'h5d == csr_addr[9:0] ? reg_csr_93 : _GEN_92; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_94 = 10'h5e == csr_addr[9:0] ? reg_csr_94 : _GEN_93; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_95 = 10'h5f == csr_addr[9:0] ? reg_csr_95 : _GEN_94; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_96 = 10'h60 == csr_addr[9:0] ? reg_csr_96 : _GEN_95; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_97 = 10'h61 == csr_addr[9:0] ? reg_csr_97 : _GEN_96; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_98 = 10'h62 == csr_addr[9:0] ? reg_csr_98 : _GEN_97; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_99 = 10'h63 == csr_addr[9:0] ? reg_csr_99 : _GEN_98; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_100 = 10'h64 == csr_addr[9:0] ? reg_csr_100 : _GEN_99; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_101 = 10'h65 == csr_addr[9:0] ? reg_csr_101 : _GEN_100; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_102 = 10'h66 == csr_addr[9:0] ? reg_csr_102 : _GEN_101; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_103 = 10'h67 == csr_addr[9:0] ? reg_csr_103 : _GEN_102; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_104 = 10'h68 == csr_addr[9:0] ? reg_csr_104 : _GEN_103; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_105 = 10'h69 == csr_addr[9:0] ? reg_csr_105 : _GEN_104; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_106 = 10'h6a == csr_addr[9:0] ? reg_csr_106 : _GEN_105; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_107 = 10'h6b == csr_addr[9:0] ? reg_csr_107 : _GEN_106; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_108 = 10'h6c == csr_addr[9:0] ? reg_csr_108 : _GEN_107; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_109 = 10'h6d == csr_addr[9:0] ? reg_csr_109 : _GEN_108; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_110 = 10'h6e == csr_addr[9:0] ? reg_csr_110 : _GEN_109; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_111 = 10'h6f == csr_addr[9:0] ? reg_csr_111 : _GEN_110; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_112 = 10'h70 == csr_addr[9:0] ? reg_csr_112 : _GEN_111; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_113 = 10'h71 == csr_addr[9:0] ? reg_csr_113 : _GEN_112; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_114 = 10'h72 == csr_addr[9:0] ? reg_csr_114 : _GEN_113; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_115 = 10'h73 == csr_addr[9:0] ? reg_csr_115 : _GEN_114; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_116 = 10'h74 == csr_addr[9:0] ? reg_csr_116 : _GEN_115; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_117 = 10'h75 == csr_addr[9:0] ? reg_csr_117 : _GEN_116; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_118 = 10'h76 == csr_addr[9:0] ? reg_csr_118 : _GEN_117; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_119 = 10'h77 == csr_addr[9:0] ? reg_csr_119 : _GEN_118; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_120 = 10'h78 == csr_addr[9:0] ? reg_csr_120 : _GEN_119; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_121 = 10'h79 == csr_addr[9:0] ? reg_csr_121 : _GEN_120; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_122 = 10'h7a == csr_addr[9:0] ? reg_csr_122 : _GEN_121; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_123 = 10'h7b == csr_addr[9:0] ? reg_csr_123 : _GEN_122; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_124 = 10'h7c == csr_addr[9:0] ? reg_csr_124 : _GEN_123; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_125 = 10'h7d == csr_addr[9:0] ? reg_csr_125 : _GEN_124; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_126 = 10'h7e == csr_addr[9:0] ? reg_csr_126 : _GEN_125; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_127 = 10'h7f == csr_addr[9:0] ? reg_csr_127 : _GEN_126; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_128 = 10'h80 == csr_addr[9:0] ? reg_csr_128 : _GEN_127; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_129 = 10'h81 == csr_addr[9:0] ? reg_csr_129 : _GEN_128; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_130 = 10'h82 == csr_addr[9:0] ? reg_csr_130 : _GEN_129; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_131 = 10'h83 == csr_addr[9:0] ? reg_csr_131 : _GEN_130; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_132 = 10'h84 == csr_addr[9:0] ? reg_csr_132 : _GEN_131; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_133 = 10'h85 == csr_addr[9:0] ? reg_csr_133 : _GEN_132; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_134 = 10'h86 == csr_addr[9:0] ? reg_csr_134 : _GEN_133; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_135 = 10'h87 == csr_addr[9:0] ? reg_csr_135 : _GEN_134; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_136 = 10'h88 == csr_addr[9:0] ? reg_csr_136 : _GEN_135; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_137 = 10'h89 == csr_addr[9:0] ? reg_csr_137 : _GEN_136; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_138 = 10'h8a == csr_addr[9:0] ? reg_csr_138 : _GEN_137; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_139 = 10'h8b == csr_addr[9:0] ? reg_csr_139 : _GEN_138; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_140 = 10'h8c == csr_addr[9:0] ? reg_csr_140 : _GEN_139; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_141 = 10'h8d == csr_addr[9:0] ? reg_csr_141 : _GEN_140; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_142 = 10'h8e == csr_addr[9:0] ? reg_csr_142 : _GEN_141; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_143 = 10'h8f == csr_addr[9:0] ? reg_csr_143 : _GEN_142; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_144 = 10'h90 == csr_addr[9:0] ? reg_csr_144 : _GEN_143; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_145 = 10'h91 == csr_addr[9:0] ? reg_csr_145 : _GEN_144; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_146 = 10'h92 == csr_addr[9:0] ? reg_csr_146 : _GEN_145; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_147 = 10'h93 == csr_addr[9:0] ? reg_csr_147 : _GEN_146; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_148 = 10'h94 == csr_addr[9:0] ? reg_csr_148 : _GEN_147; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_149 = 10'h95 == csr_addr[9:0] ? reg_csr_149 : _GEN_148; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_150 = 10'h96 == csr_addr[9:0] ? reg_csr_150 : _GEN_149; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_151 = 10'h97 == csr_addr[9:0] ? reg_csr_151 : _GEN_150; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_152 = 10'h98 == csr_addr[9:0] ? reg_csr_152 : _GEN_151; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_153 = 10'h99 == csr_addr[9:0] ? reg_csr_153 : _GEN_152; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_154 = 10'h9a == csr_addr[9:0] ? reg_csr_154 : _GEN_153; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_155 = 10'h9b == csr_addr[9:0] ? reg_csr_155 : _GEN_154; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_156 = 10'h9c == csr_addr[9:0] ? reg_csr_156 : _GEN_155; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_157 = 10'h9d == csr_addr[9:0] ? reg_csr_157 : _GEN_156; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_158 = 10'h9e == csr_addr[9:0] ? reg_csr_158 : _GEN_157; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_159 = 10'h9f == csr_addr[9:0] ? reg_csr_159 : _GEN_158; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_160 = 10'ha0 == csr_addr[9:0] ? reg_csr_160 : _GEN_159; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_161 = 10'ha1 == csr_addr[9:0] ? reg_csr_161 : _GEN_160; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_162 = 10'ha2 == csr_addr[9:0] ? reg_csr_162 : _GEN_161; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_163 = 10'ha3 == csr_addr[9:0] ? reg_csr_163 : _GEN_162; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_164 = 10'ha4 == csr_addr[9:0] ? reg_csr_164 : _GEN_163; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_165 = 10'ha5 == csr_addr[9:0] ? reg_csr_165 : _GEN_164; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_166 = 10'ha6 == csr_addr[9:0] ? reg_csr_166 : _GEN_165; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_167 = 10'ha7 == csr_addr[9:0] ? reg_csr_167 : _GEN_166; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_168 = 10'ha8 == csr_addr[9:0] ? reg_csr_168 : _GEN_167; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_169 = 10'ha9 == csr_addr[9:0] ? reg_csr_169 : _GEN_168; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_170 = 10'haa == csr_addr[9:0] ? reg_csr_170 : _GEN_169; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_171 = 10'hab == csr_addr[9:0] ? reg_csr_171 : _GEN_170; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_172 = 10'hac == csr_addr[9:0] ? reg_csr_172 : _GEN_171; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_173 = 10'had == csr_addr[9:0] ? reg_csr_173 : _GEN_172; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_174 = 10'hae == csr_addr[9:0] ? reg_csr_174 : _GEN_173; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_175 = 10'haf == csr_addr[9:0] ? reg_csr_175 : _GEN_174; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_176 = 10'hb0 == csr_addr[9:0] ? reg_csr_176 : _GEN_175; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_177 = 10'hb1 == csr_addr[9:0] ? reg_csr_177 : _GEN_176; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_178 = 10'hb2 == csr_addr[9:0] ? reg_csr_178 : _GEN_177; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_179 = 10'hb3 == csr_addr[9:0] ? reg_csr_179 : _GEN_178; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_180 = 10'hb4 == csr_addr[9:0] ? reg_csr_180 : _GEN_179; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_181 = 10'hb5 == csr_addr[9:0] ? reg_csr_181 : _GEN_180; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_182 = 10'hb6 == csr_addr[9:0] ? reg_csr_182 : _GEN_181; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_183 = 10'hb7 == csr_addr[9:0] ? reg_csr_183 : _GEN_182; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_184 = 10'hb8 == csr_addr[9:0] ? reg_csr_184 : _GEN_183; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_185 = 10'hb9 == csr_addr[9:0] ? reg_csr_185 : _GEN_184; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_186 = 10'hba == csr_addr[9:0] ? reg_csr_186 : _GEN_185; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_187 = 10'hbb == csr_addr[9:0] ? reg_csr_187 : _GEN_186; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_188 = 10'hbc == csr_addr[9:0] ? reg_csr_188 : _GEN_187; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_189 = 10'hbd == csr_addr[9:0] ? reg_csr_189 : _GEN_188; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_190 = 10'hbe == csr_addr[9:0] ? reg_csr_190 : _GEN_189; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_191 = 10'hbf == csr_addr[9:0] ? reg_csr_191 : _GEN_190; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_192 = 10'hc0 == csr_addr[9:0] ? reg_csr_192 : _GEN_191; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_193 = 10'hc1 == csr_addr[9:0] ? reg_csr_193 : _GEN_192; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_194 = 10'hc2 == csr_addr[9:0] ? reg_csr_194 : _GEN_193; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_195 = 10'hc3 == csr_addr[9:0] ? reg_csr_195 : _GEN_194; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_196 = 10'hc4 == csr_addr[9:0] ? reg_csr_196 : _GEN_195; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_197 = 10'hc5 == csr_addr[9:0] ? reg_csr_197 : _GEN_196; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_198 = 10'hc6 == csr_addr[9:0] ? reg_csr_198 : _GEN_197; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_199 = 10'hc7 == csr_addr[9:0] ? reg_csr_199 : _GEN_198; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_200 = 10'hc8 == csr_addr[9:0] ? reg_csr_200 : _GEN_199; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_201 = 10'hc9 == csr_addr[9:0] ? reg_csr_201 : _GEN_200; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_202 = 10'hca == csr_addr[9:0] ? reg_csr_202 : _GEN_201; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_203 = 10'hcb == csr_addr[9:0] ? reg_csr_203 : _GEN_202; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_204 = 10'hcc == csr_addr[9:0] ? reg_csr_204 : _GEN_203; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_205 = 10'hcd == csr_addr[9:0] ? reg_csr_205 : _GEN_204; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_206 = 10'hce == csr_addr[9:0] ? reg_csr_206 : _GEN_205; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_207 = 10'hcf == csr_addr[9:0] ? reg_csr_207 : _GEN_206; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_208 = 10'hd0 == csr_addr[9:0] ? reg_csr_208 : _GEN_207; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_209 = 10'hd1 == csr_addr[9:0] ? reg_csr_209 : _GEN_208; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_210 = 10'hd2 == csr_addr[9:0] ? reg_csr_210 : _GEN_209; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_211 = 10'hd3 == csr_addr[9:0] ? reg_csr_211 : _GEN_210; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_212 = 10'hd4 == csr_addr[9:0] ? reg_csr_212 : _GEN_211; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_213 = 10'hd5 == csr_addr[9:0] ? reg_csr_213 : _GEN_212; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_214 = 10'hd6 == csr_addr[9:0] ? reg_csr_214 : _GEN_213; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_215 = 10'hd7 == csr_addr[9:0] ? reg_csr_215 : _GEN_214; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_216 = 10'hd8 == csr_addr[9:0] ? reg_csr_216 : _GEN_215; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_217 = 10'hd9 == csr_addr[9:0] ? reg_csr_217 : _GEN_216; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_218 = 10'hda == csr_addr[9:0] ? reg_csr_218 : _GEN_217; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_219 = 10'hdb == csr_addr[9:0] ? reg_csr_219 : _GEN_218; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_220 = 10'hdc == csr_addr[9:0] ? reg_csr_220 : _GEN_219; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_221 = 10'hdd == csr_addr[9:0] ? reg_csr_221 : _GEN_220; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_222 = 10'hde == csr_addr[9:0] ? reg_csr_222 : _GEN_221; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_223 = 10'hdf == csr_addr[9:0] ? reg_csr_223 : _GEN_222; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_224 = 10'he0 == csr_addr[9:0] ? reg_csr_224 : _GEN_223; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_225 = 10'he1 == csr_addr[9:0] ? reg_csr_225 : _GEN_224; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_226 = 10'he2 == csr_addr[9:0] ? reg_csr_226 : _GEN_225; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_227 = 10'he3 == csr_addr[9:0] ? reg_csr_227 : _GEN_226; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_228 = 10'he4 == csr_addr[9:0] ? reg_csr_228 : _GEN_227; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_229 = 10'he5 == csr_addr[9:0] ? reg_csr_229 : _GEN_228; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_230 = 10'he6 == csr_addr[9:0] ? reg_csr_230 : _GEN_229; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_231 = 10'he7 == csr_addr[9:0] ? reg_csr_231 : _GEN_230; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_232 = 10'he8 == csr_addr[9:0] ? reg_csr_232 : _GEN_231; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_233 = 10'he9 == csr_addr[9:0] ? reg_csr_233 : _GEN_232; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_234 = 10'hea == csr_addr[9:0] ? reg_csr_234 : _GEN_233; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_235 = 10'heb == csr_addr[9:0] ? reg_csr_235 : _GEN_234; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_236 = 10'hec == csr_addr[9:0] ? reg_csr_236 : _GEN_235; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_237 = 10'hed == csr_addr[9:0] ? reg_csr_237 : _GEN_236; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_238 = 10'hee == csr_addr[9:0] ? reg_csr_238 : _GEN_237; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_239 = 10'hef == csr_addr[9:0] ? reg_csr_239 : _GEN_238; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_240 = 10'hf0 == csr_addr[9:0] ? reg_csr_240 : _GEN_239; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_241 = 10'hf1 == csr_addr[9:0] ? reg_csr_241 : _GEN_240; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_242 = 10'hf2 == csr_addr[9:0] ? reg_csr_242 : _GEN_241; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_243 = 10'hf3 == csr_addr[9:0] ? reg_csr_243 : _GEN_242; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_244 = 10'hf4 == csr_addr[9:0] ? reg_csr_244 : _GEN_243; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_245 = 10'hf5 == csr_addr[9:0] ? reg_csr_245 : _GEN_244; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_246 = 10'hf6 == csr_addr[9:0] ? reg_csr_246 : _GEN_245; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_247 = 10'hf7 == csr_addr[9:0] ? reg_csr_247 : _GEN_246; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_248 = 10'hf8 == csr_addr[9:0] ? reg_csr_248 : _GEN_247; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_249 = 10'hf9 == csr_addr[9:0] ? reg_csr_249 : _GEN_248; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_250 = 10'hfa == csr_addr[9:0] ? reg_csr_250 : _GEN_249; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_251 = 10'hfb == csr_addr[9:0] ? reg_csr_251 : _GEN_250; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_252 = 10'hfc == csr_addr[9:0] ? reg_csr_252 : _GEN_251; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_253 = 10'hfd == csr_addr[9:0] ? reg_csr_253 : _GEN_252; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_254 = 10'hfe == csr_addr[9:0] ? reg_csr_254 : _GEN_253; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_255 = 10'hff == csr_addr[9:0] ? reg_csr_255 : _GEN_254; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_256 = 10'h100 == csr_addr[9:0] ? reg_csr_256 : _GEN_255; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_257 = 10'h101 == csr_addr[9:0] ? reg_csr_257 : _GEN_256; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_258 = 10'h102 == csr_addr[9:0] ? reg_csr_258 : _GEN_257; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_259 = 10'h103 == csr_addr[9:0] ? reg_csr_259 : _GEN_258; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_260 = 10'h104 == csr_addr[9:0] ? reg_csr_260 : _GEN_259; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_261 = 10'h105 == csr_addr[9:0] ? reg_csr_261 : _GEN_260; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_262 = 10'h106 == csr_addr[9:0] ? reg_csr_262 : _GEN_261; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_263 = 10'h107 == csr_addr[9:0] ? reg_csr_263 : _GEN_262; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_264 = 10'h108 == csr_addr[9:0] ? reg_csr_264 : _GEN_263; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_265 = 10'h109 == csr_addr[9:0] ? reg_csr_265 : _GEN_264; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_266 = 10'h10a == csr_addr[9:0] ? reg_csr_266 : _GEN_265; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_267 = 10'h10b == csr_addr[9:0] ? reg_csr_267 : _GEN_266; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_268 = 10'h10c == csr_addr[9:0] ? reg_csr_268 : _GEN_267; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_269 = 10'h10d == csr_addr[9:0] ? reg_csr_269 : _GEN_268; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_270 = 10'h10e == csr_addr[9:0] ? reg_csr_270 : _GEN_269; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_271 = 10'h10f == csr_addr[9:0] ? reg_csr_271 : _GEN_270; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_272 = 10'h110 == csr_addr[9:0] ? reg_csr_272 : _GEN_271; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_273 = 10'h111 == csr_addr[9:0] ? reg_csr_273 : _GEN_272; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_274 = 10'h112 == csr_addr[9:0] ? reg_csr_274 : _GEN_273; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_275 = 10'h113 == csr_addr[9:0] ? reg_csr_275 : _GEN_274; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_276 = 10'h114 == csr_addr[9:0] ? reg_csr_276 : _GEN_275; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_277 = 10'h115 == csr_addr[9:0] ? reg_csr_277 : _GEN_276; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_278 = 10'h116 == csr_addr[9:0] ? reg_csr_278 : _GEN_277; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_279 = 10'h117 == csr_addr[9:0] ? reg_csr_279 : _GEN_278; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_280 = 10'h118 == csr_addr[9:0] ? reg_csr_280 : _GEN_279; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_281 = 10'h119 == csr_addr[9:0] ? reg_csr_281 : _GEN_280; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_282 = 10'h11a == csr_addr[9:0] ? reg_csr_282 : _GEN_281; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_283 = 10'h11b == csr_addr[9:0] ? reg_csr_283 : _GEN_282; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_284 = 10'h11c == csr_addr[9:0] ? reg_csr_284 : _GEN_283; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_285 = 10'h11d == csr_addr[9:0] ? reg_csr_285 : _GEN_284; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_286 = 10'h11e == csr_addr[9:0] ? reg_csr_286 : _GEN_285; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_287 = 10'h11f == csr_addr[9:0] ? reg_csr_287 : _GEN_286; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_288 = 10'h120 == csr_addr[9:0] ? reg_csr_288 : _GEN_287; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_289 = 10'h121 == csr_addr[9:0] ? reg_csr_289 : _GEN_288; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_290 = 10'h122 == csr_addr[9:0] ? reg_csr_290 : _GEN_289; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_291 = 10'h123 == csr_addr[9:0] ? reg_csr_291 : _GEN_290; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_292 = 10'h124 == csr_addr[9:0] ? reg_csr_292 : _GEN_291; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_293 = 10'h125 == csr_addr[9:0] ? reg_csr_293 : _GEN_292; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_294 = 10'h126 == csr_addr[9:0] ? reg_csr_294 : _GEN_293; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_295 = 10'h127 == csr_addr[9:0] ? reg_csr_295 : _GEN_294; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_296 = 10'h128 == csr_addr[9:0] ? reg_csr_296 : _GEN_295; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_297 = 10'h129 == csr_addr[9:0] ? reg_csr_297 : _GEN_296; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_298 = 10'h12a == csr_addr[9:0] ? reg_csr_298 : _GEN_297; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_299 = 10'h12b == csr_addr[9:0] ? reg_csr_299 : _GEN_298; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_300 = 10'h12c == csr_addr[9:0] ? reg_csr_300 : _GEN_299; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_301 = 10'h12d == csr_addr[9:0] ? reg_csr_301 : _GEN_300; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_302 = 10'h12e == csr_addr[9:0] ? reg_csr_302 : _GEN_301; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_303 = 10'h12f == csr_addr[9:0] ? reg_csr_303 : _GEN_302; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_304 = 10'h130 == csr_addr[9:0] ? reg_csr_304 : _GEN_303; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_305 = 10'h131 == csr_addr[9:0] ? reg_csr_305 : _GEN_304; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_306 = 10'h132 == csr_addr[9:0] ? reg_csr_306 : _GEN_305; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_307 = 10'h133 == csr_addr[9:0] ? reg_csr_307 : _GEN_306; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_308 = 10'h134 == csr_addr[9:0] ? reg_csr_308 : _GEN_307; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_309 = 10'h135 == csr_addr[9:0] ? reg_csr_309 : _GEN_308; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_310 = 10'h136 == csr_addr[9:0] ? reg_csr_310 : _GEN_309; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_311 = 10'h137 == csr_addr[9:0] ? reg_csr_311 : _GEN_310; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_312 = 10'h138 == csr_addr[9:0] ? reg_csr_312 : _GEN_311; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_313 = 10'h139 == csr_addr[9:0] ? reg_csr_313 : _GEN_312; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_314 = 10'h13a == csr_addr[9:0] ? reg_csr_314 : _GEN_313; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_315 = 10'h13b == csr_addr[9:0] ? reg_csr_315 : _GEN_314; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_316 = 10'h13c == csr_addr[9:0] ? reg_csr_316 : _GEN_315; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_317 = 10'h13d == csr_addr[9:0] ? reg_csr_317 : _GEN_316; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_318 = 10'h13e == csr_addr[9:0] ? reg_csr_318 : _GEN_317; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_319 = 10'h13f == csr_addr[9:0] ? reg_csr_319 : _GEN_318; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_320 = 10'h140 == csr_addr[9:0] ? reg_csr_320 : _GEN_319; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_321 = 10'h141 == csr_addr[9:0] ? reg_csr_321 : _GEN_320; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_322 = 10'h142 == csr_addr[9:0] ? reg_csr_322 : _GEN_321; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_323 = 10'h143 == csr_addr[9:0] ? reg_csr_323 : _GEN_322; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_324 = 10'h144 == csr_addr[9:0] ? reg_csr_324 : _GEN_323; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_325 = 10'h145 == csr_addr[9:0] ? reg_csr_325 : _GEN_324; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_326 = 10'h146 == csr_addr[9:0] ? reg_csr_326 : _GEN_325; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_327 = 10'h147 == csr_addr[9:0] ? reg_csr_327 : _GEN_326; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_328 = 10'h148 == csr_addr[9:0] ? reg_csr_328 : _GEN_327; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_329 = 10'h149 == csr_addr[9:0] ? reg_csr_329 : _GEN_328; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_330 = 10'h14a == csr_addr[9:0] ? reg_csr_330 : _GEN_329; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_331 = 10'h14b == csr_addr[9:0] ? reg_csr_331 : _GEN_330; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_332 = 10'h14c == csr_addr[9:0] ? reg_csr_332 : _GEN_331; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_333 = 10'h14d == csr_addr[9:0] ? reg_csr_333 : _GEN_332; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_334 = 10'h14e == csr_addr[9:0] ? reg_csr_334 : _GEN_333; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_335 = 10'h14f == csr_addr[9:0] ? reg_csr_335 : _GEN_334; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_336 = 10'h150 == csr_addr[9:0] ? reg_csr_336 : _GEN_335; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_337 = 10'h151 == csr_addr[9:0] ? reg_csr_337 : _GEN_336; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_338 = 10'h152 == csr_addr[9:0] ? reg_csr_338 : _GEN_337; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_339 = 10'h153 == csr_addr[9:0] ? reg_csr_339 : _GEN_338; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_340 = 10'h154 == csr_addr[9:0] ? reg_csr_340 : _GEN_339; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_341 = 10'h155 == csr_addr[9:0] ? reg_csr_341 : _GEN_340; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_342 = 10'h156 == csr_addr[9:0] ? reg_csr_342 : _GEN_341; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_343 = 10'h157 == csr_addr[9:0] ? reg_csr_343 : _GEN_342; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_344 = 10'h158 == csr_addr[9:0] ? reg_csr_344 : _GEN_343; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_345 = 10'h159 == csr_addr[9:0] ? reg_csr_345 : _GEN_344; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_346 = 10'h15a == csr_addr[9:0] ? reg_csr_346 : _GEN_345; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_347 = 10'h15b == csr_addr[9:0] ? reg_csr_347 : _GEN_346; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_348 = 10'h15c == csr_addr[9:0] ? reg_csr_348 : _GEN_347; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_349 = 10'h15d == csr_addr[9:0] ? reg_csr_349 : _GEN_348; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_350 = 10'h15e == csr_addr[9:0] ? reg_csr_350 : _GEN_349; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_351 = 10'h15f == csr_addr[9:0] ? reg_csr_351 : _GEN_350; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_352 = 10'h160 == csr_addr[9:0] ? reg_csr_352 : _GEN_351; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_353 = 10'h161 == csr_addr[9:0] ? reg_csr_353 : _GEN_352; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_354 = 10'h162 == csr_addr[9:0] ? reg_csr_354 : _GEN_353; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_355 = 10'h163 == csr_addr[9:0] ? reg_csr_355 : _GEN_354; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_356 = 10'h164 == csr_addr[9:0] ? reg_csr_356 : _GEN_355; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_357 = 10'h165 == csr_addr[9:0] ? reg_csr_357 : _GEN_356; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_358 = 10'h166 == csr_addr[9:0] ? reg_csr_358 : _GEN_357; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_359 = 10'h167 == csr_addr[9:0] ? reg_csr_359 : _GEN_358; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_360 = 10'h168 == csr_addr[9:0] ? reg_csr_360 : _GEN_359; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_361 = 10'h169 == csr_addr[9:0] ? reg_csr_361 : _GEN_360; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_362 = 10'h16a == csr_addr[9:0] ? reg_csr_362 : _GEN_361; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_363 = 10'h16b == csr_addr[9:0] ? reg_csr_363 : _GEN_362; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_364 = 10'h16c == csr_addr[9:0] ? reg_csr_364 : _GEN_363; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_365 = 10'h16d == csr_addr[9:0] ? reg_csr_365 : _GEN_364; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_366 = 10'h16e == csr_addr[9:0] ? reg_csr_366 : _GEN_365; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_367 = 10'h16f == csr_addr[9:0] ? reg_csr_367 : _GEN_366; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_368 = 10'h170 == csr_addr[9:0] ? reg_csr_368 : _GEN_367; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_369 = 10'h171 == csr_addr[9:0] ? reg_csr_369 : _GEN_368; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_370 = 10'h172 == csr_addr[9:0] ? reg_csr_370 : _GEN_369; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_371 = 10'h173 == csr_addr[9:0] ? reg_csr_371 : _GEN_370; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_372 = 10'h174 == csr_addr[9:0] ? reg_csr_372 : _GEN_371; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_373 = 10'h175 == csr_addr[9:0] ? reg_csr_373 : _GEN_372; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_374 = 10'h176 == csr_addr[9:0] ? reg_csr_374 : _GEN_373; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_375 = 10'h177 == csr_addr[9:0] ? reg_csr_375 : _GEN_374; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_376 = 10'h178 == csr_addr[9:0] ? reg_csr_376 : _GEN_375; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_377 = 10'h179 == csr_addr[9:0] ? reg_csr_377 : _GEN_376; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_378 = 10'h17a == csr_addr[9:0] ? reg_csr_378 : _GEN_377; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_379 = 10'h17b == csr_addr[9:0] ? reg_csr_379 : _GEN_378; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_380 = 10'h17c == csr_addr[9:0] ? reg_csr_380 : _GEN_379; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_381 = 10'h17d == csr_addr[9:0] ? reg_csr_381 : _GEN_380; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_382 = 10'h17e == csr_addr[9:0] ? reg_csr_382 : _GEN_381; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_383 = 10'h17f == csr_addr[9:0] ? reg_csr_383 : _GEN_382; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_384 = 10'h180 == csr_addr[9:0] ? reg_csr_384 : _GEN_383; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_385 = 10'h181 == csr_addr[9:0] ? reg_csr_385 : _GEN_384; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_386 = 10'h182 == csr_addr[9:0] ? reg_csr_386 : _GEN_385; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_387 = 10'h183 == csr_addr[9:0] ? reg_csr_387 : _GEN_386; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_388 = 10'h184 == csr_addr[9:0] ? reg_csr_388 : _GEN_387; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_389 = 10'h185 == csr_addr[9:0] ? reg_csr_389 : _GEN_388; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_390 = 10'h186 == csr_addr[9:0] ? reg_csr_390 : _GEN_389; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_391 = 10'h187 == csr_addr[9:0] ? reg_csr_391 : _GEN_390; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_392 = 10'h188 == csr_addr[9:0] ? reg_csr_392 : _GEN_391; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_393 = 10'h189 == csr_addr[9:0] ? reg_csr_393 : _GEN_392; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_394 = 10'h18a == csr_addr[9:0] ? reg_csr_394 : _GEN_393; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_395 = 10'h18b == csr_addr[9:0] ? reg_csr_395 : _GEN_394; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_396 = 10'h18c == csr_addr[9:0] ? reg_csr_396 : _GEN_395; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_397 = 10'h18d == csr_addr[9:0] ? reg_csr_397 : _GEN_396; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_398 = 10'h18e == csr_addr[9:0] ? reg_csr_398 : _GEN_397; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_399 = 10'h18f == csr_addr[9:0] ? reg_csr_399 : _GEN_398; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_400 = 10'h190 == csr_addr[9:0] ? reg_csr_400 : _GEN_399; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_401 = 10'h191 == csr_addr[9:0] ? reg_csr_401 : _GEN_400; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_402 = 10'h192 == csr_addr[9:0] ? reg_csr_402 : _GEN_401; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_403 = 10'h193 == csr_addr[9:0] ? reg_csr_403 : _GEN_402; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_404 = 10'h194 == csr_addr[9:0] ? reg_csr_404 : _GEN_403; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_405 = 10'h195 == csr_addr[9:0] ? reg_csr_405 : _GEN_404; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_406 = 10'h196 == csr_addr[9:0] ? reg_csr_406 : _GEN_405; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_407 = 10'h197 == csr_addr[9:0] ? reg_csr_407 : _GEN_406; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_408 = 10'h198 == csr_addr[9:0] ? reg_csr_408 : _GEN_407; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_409 = 10'h199 == csr_addr[9:0] ? reg_csr_409 : _GEN_408; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_410 = 10'h19a == csr_addr[9:0] ? reg_csr_410 : _GEN_409; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_411 = 10'h19b == csr_addr[9:0] ? reg_csr_411 : _GEN_410; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_412 = 10'h19c == csr_addr[9:0] ? reg_csr_412 : _GEN_411; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_413 = 10'h19d == csr_addr[9:0] ? reg_csr_413 : _GEN_412; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_414 = 10'h19e == csr_addr[9:0] ? reg_csr_414 : _GEN_413; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_415 = 10'h19f == csr_addr[9:0] ? reg_csr_415 : _GEN_414; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_416 = 10'h1a0 == csr_addr[9:0] ? reg_csr_416 : _GEN_415; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_417 = 10'h1a1 == csr_addr[9:0] ? reg_csr_417 : _GEN_416; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_418 = 10'h1a2 == csr_addr[9:0] ? reg_csr_418 : _GEN_417; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_419 = 10'h1a3 == csr_addr[9:0] ? reg_csr_419 : _GEN_418; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_420 = 10'h1a4 == csr_addr[9:0] ? reg_csr_420 : _GEN_419; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_421 = 10'h1a5 == csr_addr[9:0] ? reg_csr_421 : _GEN_420; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_422 = 10'h1a6 == csr_addr[9:0] ? reg_csr_422 : _GEN_421; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_423 = 10'h1a7 == csr_addr[9:0] ? reg_csr_423 : _GEN_422; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_424 = 10'h1a8 == csr_addr[9:0] ? reg_csr_424 : _GEN_423; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_425 = 10'h1a9 == csr_addr[9:0] ? reg_csr_425 : _GEN_424; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_426 = 10'h1aa == csr_addr[9:0] ? reg_csr_426 : _GEN_425; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_427 = 10'h1ab == csr_addr[9:0] ? reg_csr_427 : _GEN_426; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_428 = 10'h1ac == csr_addr[9:0] ? reg_csr_428 : _GEN_427; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_429 = 10'h1ad == csr_addr[9:0] ? reg_csr_429 : _GEN_428; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_430 = 10'h1ae == csr_addr[9:0] ? reg_csr_430 : _GEN_429; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_431 = 10'h1af == csr_addr[9:0] ? reg_csr_431 : _GEN_430; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_432 = 10'h1b0 == csr_addr[9:0] ? reg_csr_432 : _GEN_431; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_433 = 10'h1b1 == csr_addr[9:0] ? reg_csr_433 : _GEN_432; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_434 = 10'h1b2 == csr_addr[9:0] ? reg_csr_434 : _GEN_433; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_435 = 10'h1b3 == csr_addr[9:0] ? reg_csr_435 : _GEN_434; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_436 = 10'h1b4 == csr_addr[9:0] ? reg_csr_436 : _GEN_435; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_437 = 10'h1b5 == csr_addr[9:0] ? reg_csr_437 : _GEN_436; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_438 = 10'h1b6 == csr_addr[9:0] ? reg_csr_438 : _GEN_437; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_439 = 10'h1b7 == csr_addr[9:0] ? reg_csr_439 : _GEN_438; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_440 = 10'h1b8 == csr_addr[9:0] ? reg_csr_440 : _GEN_439; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_441 = 10'h1b9 == csr_addr[9:0] ? reg_csr_441 : _GEN_440; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_442 = 10'h1ba == csr_addr[9:0] ? reg_csr_442 : _GEN_441; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_443 = 10'h1bb == csr_addr[9:0] ? reg_csr_443 : _GEN_442; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_444 = 10'h1bc == csr_addr[9:0] ? reg_csr_444 : _GEN_443; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_445 = 10'h1bd == csr_addr[9:0] ? reg_csr_445 : _GEN_444; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_446 = 10'h1be == csr_addr[9:0] ? reg_csr_446 : _GEN_445; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_447 = 10'h1bf == csr_addr[9:0] ? reg_csr_447 : _GEN_446; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_448 = 10'h1c0 == csr_addr[9:0] ? reg_csr_448 : _GEN_447; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_449 = 10'h1c1 == csr_addr[9:0] ? reg_csr_449 : _GEN_448; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_450 = 10'h1c2 == csr_addr[9:0] ? reg_csr_450 : _GEN_449; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_451 = 10'h1c3 == csr_addr[9:0] ? reg_csr_451 : _GEN_450; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_452 = 10'h1c4 == csr_addr[9:0] ? reg_csr_452 : _GEN_451; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_453 = 10'h1c5 == csr_addr[9:0] ? reg_csr_453 : _GEN_452; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_454 = 10'h1c6 == csr_addr[9:0] ? reg_csr_454 : _GEN_453; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_455 = 10'h1c7 == csr_addr[9:0] ? reg_csr_455 : _GEN_454; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_456 = 10'h1c8 == csr_addr[9:0] ? reg_csr_456 : _GEN_455; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_457 = 10'h1c9 == csr_addr[9:0] ? reg_csr_457 : _GEN_456; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_458 = 10'h1ca == csr_addr[9:0] ? reg_csr_458 : _GEN_457; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_459 = 10'h1cb == csr_addr[9:0] ? reg_csr_459 : _GEN_458; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_460 = 10'h1cc == csr_addr[9:0] ? reg_csr_460 : _GEN_459; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_461 = 10'h1cd == csr_addr[9:0] ? reg_csr_461 : _GEN_460; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_462 = 10'h1ce == csr_addr[9:0] ? reg_csr_462 : _GEN_461; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_463 = 10'h1cf == csr_addr[9:0] ? reg_csr_463 : _GEN_462; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_464 = 10'h1d0 == csr_addr[9:0] ? reg_csr_464 : _GEN_463; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_465 = 10'h1d1 == csr_addr[9:0] ? reg_csr_465 : _GEN_464; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_466 = 10'h1d2 == csr_addr[9:0] ? reg_csr_466 : _GEN_465; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_467 = 10'h1d3 == csr_addr[9:0] ? reg_csr_467 : _GEN_466; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_468 = 10'h1d4 == csr_addr[9:0] ? reg_csr_468 : _GEN_467; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_469 = 10'h1d5 == csr_addr[9:0] ? reg_csr_469 : _GEN_468; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_470 = 10'h1d6 == csr_addr[9:0] ? reg_csr_470 : _GEN_469; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_471 = 10'h1d7 == csr_addr[9:0] ? reg_csr_471 : _GEN_470; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_472 = 10'h1d8 == csr_addr[9:0] ? reg_csr_472 : _GEN_471; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_473 = 10'h1d9 == csr_addr[9:0] ? reg_csr_473 : _GEN_472; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_474 = 10'h1da == csr_addr[9:0] ? reg_csr_474 : _GEN_473; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_475 = 10'h1db == csr_addr[9:0] ? reg_csr_475 : _GEN_474; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_476 = 10'h1dc == csr_addr[9:0] ? reg_csr_476 : _GEN_475; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_477 = 10'h1dd == csr_addr[9:0] ? reg_csr_477 : _GEN_476; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_478 = 10'h1de == csr_addr[9:0] ? reg_csr_478 : _GEN_477; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_479 = 10'h1df == csr_addr[9:0] ? reg_csr_479 : _GEN_478; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_480 = 10'h1e0 == csr_addr[9:0] ? reg_csr_480 : _GEN_479; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_481 = 10'h1e1 == csr_addr[9:0] ? reg_csr_481 : _GEN_480; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_482 = 10'h1e2 == csr_addr[9:0] ? reg_csr_482 : _GEN_481; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_483 = 10'h1e3 == csr_addr[9:0] ? reg_csr_483 : _GEN_482; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_484 = 10'h1e4 == csr_addr[9:0] ? reg_csr_484 : _GEN_483; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_485 = 10'h1e5 == csr_addr[9:0] ? reg_csr_485 : _GEN_484; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_486 = 10'h1e6 == csr_addr[9:0] ? reg_csr_486 : _GEN_485; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_487 = 10'h1e7 == csr_addr[9:0] ? reg_csr_487 : _GEN_486; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_488 = 10'h1e8 == csr_addr[9:0] ? reg_csr_488 : _GEN_487; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_489 = 10'h1e9 == csr_addr[9:0] ? reg_csr_489 : _GEN_488; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_490 = 10'h1ea == csr_addr[9:0] ? reg_csr_490 : _GEN_489; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_491 = 10'h1eb == csr_addr[9:0] ? reg_csr_491 : _GEN_490; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_492 = 10'h1ec == csr_addr[9:0] ? reg_csr_492 : _GEN_491; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_493 = 10'h1ed == csr_addr[9:0] ? reg_csr_493 : _GEN_492; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_494 = 10'h1ee == csr_addr[9:0] ? reg_csr_494 : _GEN_493; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_495 = 10'h1ef == csr_addr[9:0] ? reg_csr_495 : _GEN_494; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_496 = 10'h1f0 == csr_addr[9:0] ? reg_csr_496 : _GEN_495; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_497 = 10'h1f1 == csr_addr[9:0] ? reg_csr_497 : _GEN_496; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_498 = 10'h1f2 == csr_addr[9:0] ? reg_csr_498 : _GEN_497; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_499 = 10'h1f3 == csr_addr[9:0] ? reg_csr_499 : _GEN_498; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_500 = 10'h1f4 == csr_addr[9:0] ? reg_csr_500 : _GEN_499; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_501 = 10'h1f5 == csr_addr[9:0] ? reg_csr_501 : _GEN_500; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_502 = 10'h1f6 == csr_addr[9:0] ? reg_csr_502 : _GEN_501; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_503 = 10'h1f7 == csr_addr[9:0] ? reg_csr_503 : _GEN_502; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_504 = 10'h1f8 == csr_addr[9:0] ? reg_csr_504 : _GEN_503; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_505 = 10'h1f9 == csr_addr[9:0] ? reg_csr_505 : _GEN_504; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_506 = 10'h1fa == csr_addr[9:0] ? reg_csr_506 : _GEN_505; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_507 = 10'h1fb == csr_addr[9:0] ? reg_csr_507 : _GEN_506; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_508 = 10'h1fc == csr_addr[9:0] ? reg_csr_508 : _GEN_507; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_509 = 10'h1fd == csr_addr[9:0] ? reg_csr_509 : _GEN_508; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_510 = 10'h1fe == csr_addr[9:0] ? reg_csr_510 : _GEN_509; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_511 = 10'h1ff == csr_addr[9:0] ? reg_csr_511 : _GEN_510; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_512 = 10'h200 == csr_addr[9:0] ? reg_csr_512 : _GEN_511; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_513 = 10'h201 == csr_addr[9:0] ? reg_csr_513 : _GEN_512; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_514 = 10'h202 == csr_addr[9:0] ? reg_csr_514 : _GEN_513; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_515 = 10'h203 == csr_addr[9:0] ? reg_csr_515 : _GEN_514; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_516 = 10'h204 == csr_addr[9:0] ? reg_csr_516 : _GEN_515; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_517 = 10'h205 == csr_addr[9:0] ? reg_csr_517 : _GEN_516; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_518 = 10'h206 == csr_addr[9:0] ? reg_csr_518 : _GEN_517; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_519 = 10'h207 == csr_addr[9:0] ? reg_csr_519 : _GEN_518; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_520 = 10'h208 == csr_addr[9:0] ? reg_csr_520 : _GEN_519; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_521 = 10'h209 == csr_addr[9:0] ? reg_csr_521 : _GEN_520; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_522 = 10'h20a == csr_addr[9:0] ? reg_csr_522 : _GEN_521; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_523 = 10'h20b == csr_addr[9:0] ? reg_csr_523 : _GEN_522; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_524 = 10'h20c == csr_addr[9:0] ? reg_csr_524 : _GEN_523; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_525 = 10'h20d == csr_addr[9:0] ? reg_csr_525 : _GEN_524; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_526 = 10'h20e == csr_addr[9:0] ? reg_csr_526 : _GEN_525; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_527 = 10'h20f == csr_addr[9:0] ? reg_csr_527 : _GEN_526; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_528 = 10'h210 == csr_addr[9:0] ? reg_csr_528 : _GEN_527; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_529 = 10'h211 == csr_addr[9:0] ? reg_csr_529 : _GEN_528; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_530 = 10'h212 == csr_addr[9:0] ? reg_csr_530 : _GEN_529; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_531 = 10'h213 == csr_addr[9:0] ? reg_csr_531 : _GEN_530; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_532 = 10'h214 == csr_addr[9:0] ? reg_csr_532 : _GEN_531; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_533 = 10'h215 == csr_addr[9:0] ? reg_csr_533 : _GEN_532; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_534 = 10'h216 == csr_addr[9:0] ? reg_csr_534 : _GEN_533; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_535 = 10'h217 == csr_addr[9:0] ? reg_csr_535 : _GEN_534; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_536 = 10'h218 == csr_addr[9:0] ? reg_csr_536 : _GEN_535; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_537 = 10'h219 == csr_addr[9:0] ? reg_csr_537 : _GEN_536; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_538 = 10'h21a == csr_addr[9:0] ? reg_csr_538 : _GEN_537; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_539 = 10'h21b == csr_addr[9:0] ? reg_csr_539 : _GEN_538; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_540 = 10'h21c == csr_addr[9:0] ? reg_csr_540 : _GEN_539; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_541 = 10'h21d == csr_addr[9:0] ? reg_csr_541 : _GEN_540; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_542 = 10'h21e == csr_addr[9:0] ? reg_csr_542 : _GEN_541; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_543 = 10'h21f == csr_addr[9:0] ? reg_csr_543 : _GEN_542; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_544 = 10'h220 == csr_addr[9:0] ? reg_csr_544 : _GEN_543; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_545 = 10'h221 == csr_addr[9:0] ? reg_csr_545 : _GEN_544; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_546 = 10'h222 == csr_addr[9:0] ? reg_csr_546 : _GEN_545; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_547 = 10'h223 == csr_addr[9:0] ? reg_csr_547 : _GEN_546; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_548 = 10'h224 == csr_addr[9:0] ? reg_csr_548 : _GEN_547; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_549 = 10'h225 == csr_addr[9:0] ? reg_csr_549 : _GEN_548; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_550 = 10'h226 == csr_addr[9:0] ? reg_csr_550 : _GEN_549; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_551 = 10'h227 == csr_addr[9:0] ? reg_csr_551 : _GEN_550; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_552 = 10'h228 == csr_addr[9:0] ? reg_csr_552 : _GEN_551; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_553 = 10'h229 == csr_addr[9:0] ? reg_csr_553 : _GEN_552; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_554 = 10'h22a == csr_addr[9:0] ? reg_csr_554 : _GEN_553; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_555 = 10'h22b == csr_addr[9:0] ? reg_csr_555 : _GEN_554; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_556 = 10'h22c == csr_addr[9:0] ? reg_csr_556 : _GEN_555; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_557 = 10'h22d == csr_addr[9:0] ? reg_csr_557 : _GEN_556; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_558 = 10'h22e == csr_addr[9:0] ? reg_csr_558 : _GEN_557; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_559 = 10'h22f == csr_addr[9:0] ? reg_csr_559 : _GEN_558; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_560 = 10'h230 == csr_addr[9:0] ? reg_csr_560 : _GEN_559; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_561 = 10'h231 == csr_addr[9:0] ? reg_csr_561 : _GEN_560; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_562 = 10'h232 == csr_addr[9:0] ? reg_csr_562 : _GEN_561; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_563 = 10'h233 == csr_addr[9:0] ? reg_csr_563 : _GEN_562; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_564 = 10'h234 == csr_addr[9:0] ? reg_csr_564 : _GEN_563; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_565 = 10'h235 == csr_addr[9:0] ? reg_csr_565 : _GEN_564; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_566 = 10'h236 == csr_addr[9:0] ? reg_csr_566 : _GEN_565; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_567 = 10'h237 == csr_addr[9:0] ? reg_csr_567 : _GEN_566; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_568 = 10'h238 == csr_addr[9:0] ? reg_csr_568 : _GEN_567; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_569 = 10'h239 == csr_addr[9:0] ? reg_csr_569 : _GEN_568; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_570 = 10'h23a == csr_addr[9:0] ? reg_csr_570 : _GEN_569; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_571 = 10'h23b == csr_addr[9:0] ? reg_csr_571 : _GEN_570; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_572 = 10'h23c == csr_addr[9:0] ? reg_csr_572 : _GEN_571; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_573 = 10'h23d == csr_addr[9:0] ? reg_csr_573 : _GEN_572; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_574 = 10'h23e == csr_addr[9:0] ? reg_csr_574 : _GEN_573; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_575 = 10'h23f == csr_addr[9:0] ? reg_csr_575 : _GEN_574; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_576 = 10'h240 == csr_addr[9:0] ? reg_csr_576 : _GEN_575; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_577 = 10'h241 == csr_addr[9:0] ? reg_csr_577 : _GEN_576; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_578 = 10'h242 == csr_addr[9:0] ? reg_csr_578 : _GEN_577; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_579 = 10'h243 == csr_addr[9:0] ? reg_csr_579 : _GEN_578; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_580 = 10'h244 == csr_addr[9:0] ? reg_csr_580 : _GEN_579; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_581 = 10'h245 == csr_addr[9:0] ? reg_csr_581 : _GEN_580; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_582 = 10'h246 == csr_addr[9:0] ? reg_csr_582 : _GEN_581; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_583 = 10'h247 == csr_addr[9:0] ? reg_csr_583 : _GEN_582; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_584 = 10'h248 == csr_addr[9:0] ? reg_csr_584 : _GEN_583; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_585 = 10'h249 == csr_addr[9:0] ? reg_csr_585 : _GEN_584; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_586 = 10'h24a == csr_addr[9:0] ? reg_csr_586 : _GEN_585; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_587 = 10'h24b == csr_addr[9:0] ? reg_csr_587 : _GEN_586; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_588 = 10'h24c == csr_addr[9:0] ? reg_csr_588 : _GEN_587; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_589 = 10'h24d == csr_addr[9:0] ? reg_csr_589 : _GEN_588; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_590 = 10'h24e == csr_addr[9:0] ? reg_csr_590 : _GEN_589; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_591 = 10'h24f == csr_addr[9:0] ? reg_csr_591 : _GEN_590; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_592 = 10'h250 == csr_addr[9:0] ? reg_csr_592 : _GEN_591; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_593 = 10'h251 == csr_addr[9:0] ? reg_csr_593 : _GEN_592; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_594 = 10'h252 == csr_addr[9:0] ? reg_csr_594 : _GEN_593; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_595 = 10'h253 == csr_addr[9:0] ? reg_csr_595 : _GEN_594; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_596 = 10'h254 == csr_addr[9:0] ? reg_csr_596 : _GEN_595; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_597 = 10'h255 == csr_addr[9:0] ? reg_csr_597 : _GEN_596; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_598 = 10'h256 == csr_addr[9:0] ? reg_csr_598 : _GEN_597; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_599 = 10'h257 == csr_addr[9:0] ? reg_csr_599 : _GEN_598; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_600 = 10'h258 == csr_addr[9:0] ? reg_csr_600 : _GEN_599; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_601 = 10'h259 == csr_addr[9:0] ? reg_csr_601 : _GEN_600; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_602 = 10'h25a == csr_addr[9:0] ? reg_csr_602 : _GEN_601; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_603 = 10'h25b == csr_addr[9:0] ? reg_csr_603 : _GEN_602; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_604 = 10'h25c == csr_addr[9:0] ? reg_csr_604 : _GEN_603; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_605 = 10'h25d == csr_addr[9:0] ? reg_csr_605 : _GEN_604; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_606 = 10'h25e == csr_addr[9:0] ? reg_csr_606 : _GEN_605; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_607 = 10'h25f == csr_addr[9:0] ? reg_csr_607 : _GEN_606; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_608 = 10'h260 == csr_addr[9:0] ? reg_csr_608 : _GEN_607; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_609 = 10'h261 == csr_addr[9:0] ? reg_csr_609 : _GEN_608; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_610 = 10'h262 == csr_addr[9:0] ? reg_csr_610 : _GEN_609; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_611 = 10'h263 == csr_addr[9:0] ? reg_csr_611 : _GEN_610; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_612 = 10'h264 == csr_addr[9:0] ? reg_csr_612 : _GEN_611; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_613 = 10'h265 == csr_addr[9:0] ? reg_csr_613 : _GEN_612; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_614 = 10'h266 == csr_addr[9:0] ? reg_csr_614 : _GEN_613; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_615 = 10'h267 == csr_addr[9:0] ? reg_csr_615 : _GEN_614; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_616 = 10'h268 == csr_addr[9:0] ? reg_csr_616 : _GEN_615; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_617 = 10'h269 == csr_addr[9:0] ? reg_csr_617 : _GEN_616; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_618 = 10'h26a == csr_addr[9:0] ? reg_csr_618 : _GEN_617; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_619 = 10'h26b == csr_addr[9:0] ? reg_csr_619 : _GEN_618; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_620 = 10'h26c == csr_addr[9:0] ? reg_csr_620 : _GEN_619; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_621 = 10'h26d == csr_addr[9:0] ? reg_csr_621 : _GEN_620; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_622 = 10'h26e == csr_addr[9:0] ? reg_csr_622 : _GEN_621; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_623 = 10'h26f == csr_addr[9:0] ? reg_csr_623 : _GEN_622; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_624 = 10'h270 == csr_addr[9:0] ? reg_csr_624 : _GEN_623; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_625 = 10'h271 == csr_addr[9:0] ? reg_csr_625 : _GEN_624; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_626 = 10'h272 == csr_addr[9:0] ? reg_csr_626 : _GEN_625; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_627 = 10'h273 == csr_addr[9:0] ? reg_csr_627 : _GEN_626; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_628 = 10'h274 == csr_addr[9:0] ? reg_csr_628 : _GEN_627; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_629 = 10'h275 == csr_addr[9:0] ? reg_csr_629 : _GEN_628; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_630 = 10'h276 == csr_addr[9:0] ? reg_csr_630 : _GEN_629; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_631 = 10'h277 == csr_addr[9:0] ? reg_csr_631 : _GEN_630; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_632 = 10'h278 == csr_addr[9:0] ? reg_csr_632 : _GEN_631; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_633 = 10'h279 == csr_addr[9:0] ? reg_csr_633 : _GEN_632; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_634 = 10'h27a == csr_addr[9:0] ? reg_csr_634 : _GEN_633; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_635 = 10'h27b == csr_addr[9:0] ? reg_csr_635 : _GEN_634; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_636 = 10'h27c == csr_addr[9:0] ? reg_csr_636 : _GEN_635; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_637 = 10'h27d == csr_addr[9:0] ? reg_csr_637 : _GEN_636; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_638 = 10'h27e == csr_addr[9:0] ? reg_csr_638 : _GEN_637; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_639 = 10'h27f == csr_addr[9:0] ? reg_csr_639 : _GEN_638; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_640 = 10'h280 == csr_addr[9:0] ? reg_csr_640 : _GEN_639; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_641 = 10'h281 == csr_addr[9:0] ? reg_csr_641 : _GEN_640; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_642 = 10'h282 == csr_addr[9:0] ? reg_csr_642 : _GEN_641; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_643 = 10'h283 == csr_addr[9:0] ? reg_csr_643 : _GEN_642; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_644 = 10'h284 == csr_addr[9:0] ? reg_csr_644 : _GEN_643; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_645 = 10'h285 == csr_addr[9:0] ? reg_csr_645 : _GEN_644; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_646 = 10'h286 == csr_addr[9:0] ? reg_csr_646 : _GEN_645; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_647 = 10'h287 == csr_addr[9:0] ? reg_csr_647 : _GEN_646; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_648 = 10'h288 == csr_addr[9:0] ? reg_csr_648 : _GEN_647; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_649 = 10'h289 == csr_addr[9:0] ? reg_csr_649 : _GEN_648; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_650 = 10'h28a == csr_addr[9:0] ? reg_csr_650 : _GEN_649; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_651 = 10'h28b == csr_addr[9:0] ? reg_csr_651 : _GEN_650; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_652 = 10'h28c == csr_addr[9:0] ? reg_csr_652 : _GEN_651; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_653 = 10'h28d == csr_addr[9:0] ? reg_csr_653 : _GEN_652; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_654 = 10'h28e == csr_addr[9:0] ? reg_csr_654 : _GEN_653; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_655 = 10'h28f == csr_addr[9:0] ? reg_csr_655 : _GEN_654; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_656 = 10'h290 == csr_addr[9:0] ? reg_csr_656 : _GEN_655; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_657 = 10'h291 == csr_addr[9:0] ? reg_csr_657 : _GEN_656; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_658 = 10'h292 == csr_addr[9:0] ? reg_csr_658 : _GEN_657; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_659 = 10'h293 == csr_addr[9:0] ? reg_csr_659 : _GEN_658; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_660 = 10'h294 == csr_addr[9:0] ? reg_csr_660 : _GEN_659; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_661 = 10'h295 == csr_addr[9:0] ? reg_csr_661 : _GEN_660; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_662 = 10'h296 == csr_addr[9:0] ? reg_csr_662 : _GEN_661; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_663 = 10'h297 == csr_addr[9:0] ? reg_csr_663 : _GEN_662; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_664 = 10'h298 == csr_addr[9:0] ? reg_csr_664 : _GEN_663; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_665 = 10'h299 == csr_addr[9:0] ? reg_csr_665 : _GEN_664; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_666 = 10'h29a == csr_addr[9:0] ? reg_csr_666 : _GEN_665; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_667 = 10'h29b == csr_addr[9:0] ? reg_csr_667 : _GEN_666; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_668 = 10'h29c == csr_addr[9:0] ? reg_csr_668 : _GEN_667; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_669 = 10'h29d == csr_addr[9:0] ? reg_csr_669 : _GEN_668; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_670 = 10'h29e == csr_addr[9:0] ? reg_csr_670 : _GEN_669; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_671 = 10'h29f == csr_addr[9:0] ? reg_csr_671 : _GEN_670; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_672 = 10'h2a0 == csr_addr[9:0] ? reg_csr_672 : _GEN_671; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_673 = 10'h2a1 == csr_addr[9:0] ? reg_csr_673 : _GEN_672; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_674 = 10'h2a2 == csr_addr[9:0] ? reg_csr_674 : _GEN_673; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_675 = 10'h2a3 == csr_addr[9:0] ? reg_csr_675 : _GEN_674; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_676 = 10'h2a4 == csr_addr[9:0] ? reg_csr_676 : _GEN_675; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_677 = 10'h2a5 == csr_addr[9:0] ? reg_csr_677 : _GEN_676; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_678 = 10'h2a6 == csr_addr[9:0] ? reg_csr_678 : _GEN_677; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_679 = 10'h2a7 == csr_addr[9:0] ? reg_csr_679 : _GEN_678; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_680 = 10'h2a8 == csr_addr[9:0] ? reg_csr_680 : _GEN_679; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_681 = 10'h2a9 == csr_addr[9:0] ? reg_csr_681 : _GEN_680; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_682 = 10'h2aa == csr_addr[9:0] ? reg_csr_682 : _GEN_681; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_683 = 10'h2ab == csr_addr[9:0] ? reg_csr_683 : _GEN_682; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_684 = 10'h2ac == csr_addr[9:0] ? reg_csr_684 : _GEN_683; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_685 = 10'h2ad == csr_addr[9:0] ? reg_csr_685 : _GEN_684; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_686 = 10'h2ae == csr_addr[9:0] ? reg_csr_686 : _GEN_685; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_687 = 10'h2af == csr_addr[9:0] ? reg_csr_687 : _GEN_686; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_688 = 10'h2b0 == csr_addr[9:0] ? reg_csr_688 : _GEN_687; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_689 = 10'h2b1 == csr_addr[9:0] ? reg_csr_689 : _GEN_688; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_690 = 10'h2b2 == csr_addr[9:0] ? reg_csr_690 : _GEN_689; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_691 = 10'h2b3 == csr_addr[9:0] ? reg_csr_691 : _GEN_690; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_692 = 10'h2b4 == csr_addr[9:0] ? reg_csr_692 : _GEN_691; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_693 = 10'h2b5 == csr_addr[9:0] ? reg_csr_693 : _GEN_692; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_694 = 10'h2b6 == csr_addr[9:0] ? reg_csr_694 : _GEN_693; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_695 = 10'h2b7 == csr_addr[9:0] ? reg_csr_695 : _GEN_694; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_696 = 10'h2b8 == csr_addr[9:0] ? reg_csr_696 : _GEN_695; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_697 = 10'h2b9 == csr_addr[9:0] ? reg_csr_697 : _GEN_696; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_698 = 10'h2ba == csr_addr[9:0] ? reg_csr_698 : _GEN_697; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_699 = 10'h2bb == csr_addr[9:0] ? reg_csr_699 : _GEN_698; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_700 = 10'h2bc == csr_addr[9:0] ? reg_csr_700 : _GEN_699; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_701 = 10'h2bd == csr_addr[9:0] ? reg_csr_701 : _GEN_700; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_702 = 10'h2be == csr_addr[9:0] ? reg_csr_702 : _GEN_701; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_703 = 10'h2bf == csr_addr[9:0] ? reg_csr_703 : _GEN_702; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_704 = 10'h2c0 == csr_addr[9:0] ? reg_csr_704 : _GEN_703; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_705 = 10'h2c1 == csr_addr[9:0] ? reg_csr_705 : _GEN_704; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_706 = 10'h2c2 == csr_addr[9:0] ? reg_csr_706 : _GEN_705; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_707 = 10'h2c3 == csr_addr[9:0] ? reg_csr_707 : _GEN_706; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_708 = 10'h2c4 == csr_addr[9:0] ? reg_csr_708 : _GEN_707; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_709 = 10'h2c5 == csr_addr[9:0] ? reg_csr_709 : _GEN_708; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_710 = 10'h2c6 == csr_addr[9:0] ? reg_csr_710 : _GEN_709; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_711 = 10'h2c7 == csr_addr[9:0] ? reg_csr_711 : _GEN_710; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_712 = 10'h2c8 == csr_addr[9:0] ? reg_csr_712 : _GEN_711; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_713 = 10'h2c9 == csr_addr[9:0] ? reg_csr_713 : _GEN_712; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_714 = 10'h2ca == csr_addr[9:0] ? reg_csr_714 : _GEN_713; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_715 = 10'h2cb == csr_addr[9:0] ? reg_csr_715 : _GEN_714; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_716 = 10'h2cc == csr_addr[9:0] ? reg_csr_716 : _GEN_715; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_717 = 10'h2cd == csr_addr[9:0] ? reg_csr_717 : _GEN_716; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_718 = 10'h2ce == csr_addr[9:0] ? reg_csr_718 : _GEN_717; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_719 = 10'h2cf == csr_addr[9:0] ? reg_csr_719 : _GEN_718; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_720 = 10'h2d0 == csr_addr[9:0] ? reg_csr_720 : _GEN_719; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_721 = 10'h2d1 == csr_addr[9:0] ? reg_csr_721 : _GEN_720; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_722 = 10'h2d2 == csr_addr[9:0] ? reg_csr_722 : _GEN_721; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_723 = 10'h2d3 == csr_addr[9:0] ? reg_csr_723 : _GEN_722; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_724 = 10'h2d4 == csr_addr[9:0] ? reg_csr_724 : _GEN_723; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_725 = 10'h2d5 == csr_addr[9:0] ? reg_csr_725 : _GEN_724; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_726 = 10'h2d6 == csr_addr[9:0] ? reg_csr_726 : _GEN_725; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_727 = 10'h2d7 == csr_addr[9:0] ? reg_csr_727 : _GEN_726; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_728 = 10'h2d8 == csr_addr[9:0] ? reg_csr_728 : _GEN_727; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_729 = 10'h2d9 == csr_addr[9:0] ? reg_csr_729 : _GEN_728; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_730 = 10'h2da == csr_addr[9:0] ? reg_csr_730 : _GEN_729; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_731 = 10'h2db == csr_addr[9:0] ? reg_csr_731 : _GEN_730; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_732 = 10'h2dc == csr_addr[9:0] ? reg_csr_732 : _GEN_731; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_733 = 10'h2dd == csr_addr[9:0] ? reg_csr_733 : _GEN_732; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_734 = 10'h2de == csr_addr[9:0] ? reg_csr_734 : _GEN_733; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_735 = 10'h2df == csr_addr[9:0] ? reg_csr_735 : _GEN_734; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_736 = 10'h2e0 == csr_addr[9:0] ? reg_csr_736 : _GEN_735; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_737 = 10'h2e1 == csr_addr[9:0] ? reg_csr_737 : _GEN_736; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_738 = 10'h2e2 == csr_addr[9:0] ? reg_csr_738 : _GEN_737; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_739 = 10'h2e3 == csr_addr[9:0] ? reg_csr_739 : _GEN_738; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_740 = 10'h2e4 == csr_addr[9:0] ? reg_csr_740 : _GEN_739; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_741 = 10'h2e5 == csr_addr[9:0] ? reg_csr_741 : _GEN_740; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_742 = 10'h2e6 == csr_addr[9:0] ? reg_csr_742 : _GEN_741; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_743 = 10'h2e7 == csr_addr[9:0] ? reg_csr_743 : _GEN_742; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_744 = 10'h2e8 == csr_addr[9:0] ? reg_csr_744 : _GEN_743; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_745 = 10'h2e9 == csr_addr[9:0] ? reg_csr_745 : _GEN_744; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_746 = 10'h2ea == csr_addr[9:0] ? reg_csr_746 : _GEN_745; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_747 = 10'h2eb == csr_addr[9:0] ? reg_csr_747 : _GEN_746; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_748 = 10'h2ec == csr_addr[9:0] ? reg_csr_748 : _GEN_747; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_749 = 10'h2ed == csr_addr[9:0] ? reg_csr_749 : _GEN_748; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_750 = 10'h2ee == csr_addr[9:0] ? reg_csr_750 : _GEN_749; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_751 = 10'h2ef == csr_addr[9:0] ? reg_csr_751 : _GEN_750; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_752 = 10'h2f0 == csr_addr[9:0] ? reg_csr_752 : _GEN_751; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_753 = 10'h2f1 == csr_addr[9:0] ? reg_csr_753 : _GEN_752; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_754 = 10'h2f2 == csr_addr[9:0] ? reg_csr_754 : _GEN_753; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_755 = 10'h2f3 == csr_addr[9:0] ? reg_csr_755 : _GEN_754; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_756 = 10'h2f4 == csr_addr[9:0] ? reg_csr_756 : _GEN_755; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_757 = 10'h2f5 == csr_addr[9:0] ? reg_csr_757 : _GEN_756; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_758 = 10'h2f6 == csr_addr[9:0] ? reg_csr_758 : _GEN_757; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_759 = 10'h2f7 == csr_addr[9:0] ? reg_csr_759 : _GEN_758; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_760 = 10'h2f8 == csr_addr[9:0] ? reg_csr_760 : _GEN_759; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_761 = 10'h2f9 == csr_addr[9:0] ? reg_csr_761 : _GEN_760; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_762 = 10'h2fa == csr_addr[9:0] ? reg_csr_762 : _GEN_761; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_763 = 10'h2fb == csr_addr[9:0] ? reg_csr_763 : _GEN_762; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_764 = 10'h2fc == csr_addr[9:0] ? reg_csr_764 : _GEN_763; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_765 = 10'h2fd == csr_addr[9:0] ? reg_csr_765 : _GEN_764; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_766 = 10'h2fe == csr_addr[9:0] ? reg_csr_766 : _GEN_765; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_767 = 10'h2ff == csr_addr[9:0] ? reg_csr_767 : _GEN_766; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_768 = 10'h300 == csr_addr[9:0] ? reg_csr_768 : _GEN_767; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_769 = 10'h301 == csr_addr[9:0] ? reg_csr_769 : _GEN_768; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_770 = 10'h302 == csr_addr[9:0] ? reg_csr_770 : _GEN_769; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_771 = 10'h303 == csr_addr[9:0] ? reg_csr_771 : _GEN_770; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_772 = 10'h304 == csr_addr[9:0] ? reg_csr_772 : _GEN_771; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_773 = 10'h305 == csr_addr[9:0] ? reg_csr_773 : _GEN_772; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_774 = 10'h306 == csr_addr[9:0] ? reg_csr_774 : _GEN_773; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_775 = 10'h307 == csr_addr[9:0] ? reg_csr_775 : _GEN_774; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_776 = 10'h308 == csr_addr[9:0] ? reg_csr_776 : _GEN_775; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_777 = 10'h309 == csr_addr[9:0] ? reg_csr_777 : _GEN_776; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_778 = 10'h30a == csr_addr[9:0] ? reg_csr_778 : _GEN_777; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_779 = 10'h30b == csr_addr[9:0] ? reg_csr_779 : _GEN_778; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_780 = 10'h30c == csr_addr[9:0] ? reg_csr_780 : _GEN_779; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_781 = 10'h30d == csr_addr[9:0] ? reg_csr_781 : _GEN_780; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_782 = 10'h30e == csr_addr[9:0] ? reg_csr_782 : _GEN_781; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_783 = 10'h30f == csr_addr[9:0] ? reg_csr_783 : _GEN_782; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_784 = 10'h310 == csr_addr[9:0] ? reg_csr_784 : _GEN_783; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_785 = 10'h311 == csr_addr[9:0] ? reg_csr_785 : _GEN_784; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_786 = 10'h312 == csr_addr[9:0] ? reg_csr_786 : _GEN_785; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_787 = 10'h313 == csr_addr[9:0] ? reg_csr_787 : _GEN_786; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_788 = 10'h314 == csr_addr[9:0] ? reg_csr_788 : _GEN_787; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_789 = 10'h315 == csr_addr[9:0] ? reg_csr_789 : _GEN_788; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_790 = 10'h316 == csr_addr[9:0] ? reg_csr_790 : _GEN_789; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_791 = 10'h317 == csr_addr[9:0] ? reg_csr_791 : _GEN_790; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_792 = 10'h318 == csr_addr[9:0] ? reg_csr_792 : _GEN_791; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_793 = 10'h319 == csr_addr[9:0] ? reg_csr_793 : _GEN_792; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_794 = 10'h31a == csr_addr[9:0] ? reg_csr_794 : _GEN_793; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_795 = 10'h31b == csr_addr[9:0] ? reg_csr_795 : _GEN_794; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_796 = 10'h31c == csr_addr[9:0] ? reg_csr_796 : _GEN_795; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_797 = 10'h31d == csr_addr[9:0] ? reg_csr_797 : _GEN_796; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_798 = 10'h31e == csr_addr[9:0] ? reg_csr_798 : _GEN_797; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_799 = 10'h31f == csr_addr[9:0] ? reg_csr_799 : _GEN_798; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_800 = 10'h320 == csr_addr[9:0] ? reg_csr_800 : _GEN_799; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_801 = 10'h321 == csr_addr[9:0] ? reg_csr_801 : _GEN_800; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_802 = 10'h322 == csr_addr[9:0] ? reg_csr_802 : _GEN_801; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_803 = 10'h323 == csr_addr[9:0] ? reg_csr_803 : _GEN_802; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_804 = 10'h324 == csr_addr[9:0] ? reg_csr_804 : _GEN_803; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_805 = 10'h325 == csr_addr[9:0] ? reg_csr_805 : _GEN_804; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_806 = 10'h326 == csr_addr[9:0] ? reg_csr_806 : _GEN_805; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_807 = 10'h327 == csr_addr[9:0] ? reg_csr_807 : _GEN_806; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_808 = 10'h328 == csr_addr[9:0] ? reg_csr_808 : _GEN_807; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_809 = 10'h329 == csr_addr[9:0] ? reg_csr_809 : _GEN_808; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_810 = 10'h32a == csr_addr[9:0] ? reg_csr_810 : _GEN_809; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_811 = 10'h32b == csr_addr[9:0] ? reg_csr_811 : _GEN_810; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_812 = 10'h32c == csr_addr[9:0] ? reg_csr_812 : _GEN_811; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_813 = 10'h32d == csr_addr[9:0] ? reg_csr_813 : _GEN_812; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_814 = 10'h32e == csr_addr[9:0] ? reg_csr_814 : _GEN_813; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_815 = 10'h32f == csr_addr[9:0] ? reg_csr_815 : _GEN_814; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_816 = 10'h330 == csr_addr[9:0] ? reg_csr_816 : _GEN_815; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_817 = 10'h331 == csr_addr[9:0] ? reg_csr_817 : _GEN_816; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_818 = 10'h332 == csr_addr[9:0] ? reg_csr_818 : _GEN_817; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_819 = 10'h333 == csr_addr[9:0] ? reg_csr_819 : _GEN_818; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_820 = 10'h334 == csr_addr[9:0] ? reg_csr_820 : _GEN_819; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_821 = 10'h335 == csr_addr[9:0] ? reg_csr_821 : _GEN_820; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_822 = 10'h336 == csr_addr[9:0] ? reg_csr_822 : _GEN_821; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_823 = 10'h337 == csr_addr[9:0] ? reg_csr_823 : _GEN_822; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_824 = 10'h338 == csr_addr[9:0] ? reg_csr_824 : _GEN_823; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_825 = 10'h339 == csr_addr[9:0] ? reg_csr_825 : _GEN_824; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_826 = 10'h33a == csr_addr[9:0] ? reg_csr_826 : _GEN_825; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_827 = 10'h33b == csr_addr[9:0] ? reg_csr_827 : _GEN_826; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_828 = 10'h33c == csr_addr[9:0] ? reg_csr_828 : _GEN_827; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_829 = 10'h33d == csr_addr[9:0] ? reg_csr_829 : _GEN_828; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_830 = 10'h33e == csr_addr[9:0] ? reg_csr_830 : _GEN_829; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_831 = 10'h33f == csr_addr[9:0] ? reg_csr_831 : _GEN_830; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_832 = 10'h340 == csr_addr[9:0] ? reg_csr_832 : _GEN_831; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_833 = 10'h341 == csr_addr[9:0] ? reg_csr_833 : _GEN_832; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_834 = 10'h342 == csr_addr[9:0] ? reg_csr_834 : _GEN_833; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_835 = 10'h343 == csr_addr[9:0] ? reg_csr_835 : _GEN_834; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_836 = 10'h344 == csr_addr[9:0] ? reg_csr_836 : _GEN_835; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_837 = 10'h345 == csr_addr[9:0] ? reg_csr_837 : _GEN_836; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_838 = 10'h346 == csr_addr[9:0] ? reg_csr_838 : _GEN_837; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_839 = 10'h347 == csr_addr[9:0] ? reg_csr_839 : _GEN_838; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_840 = 10'h348 == csr_addr[9:0] ? reg_csr_840 : _GEN_839; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_841 = 10'h349 == csr_addr[9:0] ? reg_csr_841 : _GEN_840; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_842 = 10'h34a == csr_addr[9:0] ? reg_csr_842 : _GEN_841; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_843 = 10'h34b == csr_addr[9:0] ? reg_csr_843 : _GEN_842; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_844 = 10'h34c == csr_addr[9:0] ? reg_csr_844 : _GEN_843; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_845 = 10'h34d == csr_addr[9:0] ? reg_csr_845 : _GEN_844; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_846 = 10'h34e == csr_addr[9:0] ? reg_csr_846 : _GEN_845; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_847 = 10'h34f == csr_addr[9:0] ? reg_csr_847 : _GEN_846; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_848 = 10'h350 == csr_addr[9:0] ? reg_csr_848 : _GEN_847; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_849 = 10'h351 == csr_addr[9:0] ? reg_csr_849 : _GEN_848; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_850 = 10'h352 == csr_addr[9:0] ? reg_csr_850 : _GEN_849; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_851 = 10'h353 == csr_addr[9:0] ? reg_csr_851 : _GEN_850; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_852 = 10'h354 == csr_addr[9:0] ? reg_csr_852 : _GEN_851; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_853 = 10'h355 == csr_addr[9:0] ? reg_csr_853 : _GEN_852; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_854 = 10'h356 == csr_addr[9:0] ? reg_csr_854 : _GEN_853; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_855 = 10'h357 == csr_addr[9:0] ? reg_csr_855 : _GEN_854; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_856 = 10'h358 == csr_addr[9:0] ? reg_csr_856 : _GEN_855; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_857 = 10'h359 == csr_addr[9:0] ? reg_csr_857 : _GEN_856; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_858 = 10'h35a == csr_addr[9:0] ? reg_csr_858 : _GEN_857; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_859 = 10'h35b == csr_addr[9:0] ? reg_csr_859 : _GEN_858; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_860 = 10'h35c == csr_addr[9:0] ? reg_csr_860 : _GEN_859; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_861 = 10'h35d == csr_addr[9:0] ? reg_csr_861 : _GEN_860; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_862 = 10'h35e == csr_addr[9:0] ? reg_csr_862 : _GEN_861; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_863 = 10'h35f == csr_addr[9:0] ? reg_csr_863 : _GEN_862; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_864 = 10'h360 == csr_addr[9:0] ? reg_csr_864 : _GEN_863; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_865 = 10'h361 == csr_addr[9:0] ? reg_csr_865 : _GEN_864; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_866 = 10'h362 == csr_addr[9:0] ? reg_csr_866 : _GEN_865; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_867 = 10'h363 == csr_addr[9:0] ? reg_csr_867 : _GEN_866; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_868 = 10'h364 == csr_addr[9:0] ? reg_csr_868 : _GEN_867; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_869 = 10'h365 == csr_addr[9:0] ? reg_csr_869 : _GEN_868; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_870 = 10'h366 == csr_addr[9:0] ? reg_csr_870 : _GEN_869; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_871 = 10'h367 == csr_addr[9:0] ? reg_csr_871 : _GEN_870; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_872 = 10'h368 == csr_addr[9:0] ? reg_csr_872 : _GEN_871; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_873 = 10'h369 == csr_addr[9:0] ? reg_csr_873 : _GEN_872; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_874 = 10'h36a == csr_addr[9:0] ? reg_csr_874 : _GEN_873; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_875 = 10'h36b == csr_addr[9:0] ? reg_csr_875 : _GEN_874; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_876 = 10'h36c == csr_addr[9:0] ? reg_csr_876 : _GEN_875; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_877 = 10'h36d == csr_addr[9:0] ? reg_csr_877 : _GEN_876; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_878 = 10'h36e == csr_addr[9:0] ? reg_csr_878 : _GEN_877; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_879 = 10'h36f == csr_addr[9:0] ? reg_csr_879 : _GEN_878; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_880 = 10'h370 == csr_addr[9:0] ? reg_csr_880 : _GEN_879; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_881 = 10'h371 == csr_addr[9:0] ? reg_csr_881 : _GEN_880; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_882 = 10'h372 == csr_addr[9:0] ? reg_csr_882 : _GEN_881; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_883 = 10'h373 == csr_addr[9:0] ? reg_csr_883 : _GEN_882; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_884 = 10'h374 == csr_addr[9:0] ? reg_csr_884 : _GEN_883; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_885 = 10'h375 == csr_addr[9:0] ? reg_csr_885 : _GEN_884; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_886 = 10'h376 == csr_addr[9:0] ? reg_csr_886 : _GEN_885; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_887 = 10'h377 == csr_addr[9:0] ? reg_csr_887 : _GEN_886; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_888 = 10'h378 == csr_addr[9:0] ? reg_csr_888 : _GEN_887; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_889 = 10'h379 == csr_addr[9:0] ? reg_csr_889 : _GEN_888; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_890 = 10'h37a == csr_addr[9:0] ? reg_csr_890 : _GEN_889; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_891 = 10'h37b == csr_addr[9:0] ? reg_csr_891 : _GEN_890; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_892 = 10'h37c == csr_addr[9:0] ? reg_csr_892 : _GEN_891; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_893 = 10'h37d == csr_addr[9:0] ? reg_csr_893 : _GEN_892; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_894 = 10'h37e == csr_addr[9:0] ? reg_csr_894 : _GEN_893; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_895 = 10'h37f == csr_addr[9:0] ? reg_csr_895 : _GEN_894; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_896 = 10'h380 == csr_addr[9:0] ? reg_csr_896 : _GEN_895; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_897 = 10'h381 == csr_addr[9:0] ? reg_csr_897 : _GEN_896; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_898 = 10'h382 == csr_addr[9:0] ? reg_csr_898 : _GEN_897; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_899 = 10'h383 == csr_addr[9:0] ? reg_csr_899 : _GEN_898; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_900 = 10'h384 == csr_addr[9:0] ? reg_csr_900 : _GEN_899; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_901 = 10'h385 == csr_addr[9:0] ? reg_csr_901 : _GEN_900; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_902 = 10'h386 == csr_addr[9:0] ? reg_csr_902 : _GEN_901; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_903 = 10'h387 == csr_addr[9:0] ? reg_csr_903 : _GEN_902; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_904 = 10'h388 == csr_addr[9:0] ? reg_csr_904 : _GEN_903; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_905 = 10'h389 == csr_addr[9:0] ? reg_csr_905 : _GEN_904; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_906 = 10'h38a == csr_addr[9:0] ? reg_csr_906 : _GEN_905; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_907 = 10'h38b == csr_addr[9:0] ? reg_csr_907 : _GEN_906; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_908 = 10'h38c == csr_addr[9:0] ? reg_csr_908 : _GEN_907; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_909 = 10'h38d == csr_addr[9:0] ? reg_csr_909 : _GEN_908; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_910 = 10'h38e == csr_addr[9:0] ? reg_csr_910 : _GEN_909; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_911 = 10'h38f == csr_addr[9:0] ? reg_csr_911 : _GEN_910; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_912 = 10'h390 == csr_addr[9:0] ? reg_csr_912 : _GEN_911; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_913 = 10'h391 == csr_addr[9:0] ? reg_csr_913 : _GEN_912; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_914 = 10'h392 == csr_addr[9:0] ? reg_csr_914 : _GEN_913; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_915 = 10'h393 == csr_addr[9:0] ? reg_csr_915 : _GEN_914; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_916 = 10'h394 == csr_addr[9:0] ? reg_csr_916 : _GEN_915; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_917 = 10'h395 == csr_addr[9:0] ? reg_csr_917 : _GEN_916; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_918 = 10'h396 == csr_addr[9:0] ? reg_csr_918 : _GEN_917; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_919 = 10'h397 == csr_addr[9:0] ? reg_csr_919 : _GEN_918; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_920 = 10'h398 == csr_addr[9:0] ? reg_csr_920 : _GEN_919; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_921 = 10'h399 == csr_addr[9:0] ? reg_csr_921 : _GEN_920; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_922 = 10'h39a == csr_addr[9:0] ? reg_csr_922 : _GEN_921; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_923 = 10'h39b == csr_addr[9:0] ? reg_csr_923 : _GEN_922; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_924 = 10'h39c == csr_addr[9:0] ? reg_csr_924 : _GEN_923; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_925 = 10'h39d == csr_addr[9:0] ? reg_csr_925 : _GEN_924; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_926 = 10'h39e == csr_addr[9:0] ? reg_csr_926 : _GEN_925; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_927 = 10'h39f == csr_addr[9:0] ? reg_csr_927 : _GEN_926; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_928 = 10'h3a0 == csr_addr[9:0] ? reg_csr_928 : _GEN_927; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_929 = 10'h3a1 == csr_addr[9:0] ? reg_csr_929 : _GEN_928; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_930 = 10'h3a2 == csr_addr[9:0] ? reg_csr_930 : _GEN_929; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_931 = 10'h3a3 == csr_addr[9:0] ? reg_csr_931 : _GEN_930; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_932 = 10'h3a4 == csr_addr[9:0] ? reg_csr_932 : _GEN_931; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_933 = 10'h3a5 == csr_addr[9:0] ? reg_csr_933 : _GEN_932; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_934 = 10'h3a6 == csr_addr[9:0] ? reg_csr_934 : _GEN_933; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_935 = 10'h3a7 == csr_addr[9:0] ? reg_csr_935 : _GEN_934; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_936 = 10'h3a8 == csr_addr[9:0] ? reg_csr_936 : _GEN_935; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_937 = 10'h3a9 == csr_addr[9:0] ? reg_csr_937 : _GEN_936; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_938 = 10'h3aa == csr_addr[9:0] ? reg_csr_938 : _GEN_937; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_939 = 10'h3ab == csr_addr[9:0] ? reg_csr_939 : _GEN_938; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_940 = 10'h3ac == csr_addr[9:0] ? reg_csr_940 : _GEN_939; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_941 = 10'h3ad == csr_addr[9:0] ? reg_csr_941 : _GEN_940; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_942 = 10'h3ae == csr_addr[9:0] ? reg_csr_942 : _GEN_941; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_943 = 10'h3af == csr_addr[9:0] ? reg_csr_943 : _GEN_942; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_944 = 10'h3b0 == csr_addr[9:0] ? reg_csr_944 : _GEN_943; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_945 = 10'h3b1 == csr_addr[9:0] ? reg_csr_945 : _GEN_944; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_946 = 10'h3b2 == csr_addr[9:0] ? reg_csr_946 : _GEN_945; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_947 = 10'h3b3 == csr_addr[9:0] ? reg_csr_947 : _GEN_946; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_948 = 10'h3b4 == csr_addr[9:0] ? reg_csr_948 : _GEN_947; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_949 = 10'h3b5 == csr_addr[9:0] ? reg_csr_949 : _GEN_948; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_950 = 10'h3b6 == csr_addr[9:0] ? reg_csr_950 : _GEN_949; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_951 = 10'h3b7 == csr_addr[9:0] ? reg_csr_951 : _GEN_950; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_952 = 10'h3b8 == csr_addr[9:0] ? reg_csr_952 : _GEN_951; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_953 = 10'h3b9 == csr_addr[9:0] ? reg_csr_953 : _GEN_952; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_954 = 10'h3ba == csr_addr[9:0] ? reg_csr_954 : _GEN_953; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_955 = 10'h3bb == csr_addr[9:0] ? reg_csr_955 : _GEN_954; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_956 = 10'h3bc == csr_addr[9:0] ? reg_csr_956 : _GEN_955; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_957 = 10'h3bd == csr_addr[9:0] ? reg_csr_957 : _GEN_956; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_958 = 10'h3be == csr_addr[9:0] ? reg_csr_958 : _GEN_957; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_959 = 10'h3bf == csr_addr[9:0] ? reg_csr_959 : _GEN_958; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_960 = 10'h3c0 == csr_addr[9:0] ? reg_csr_960 : _GEN_959; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_961 = 10'h3c1 == csr_addr[9:0] ? reg_csr_961 : _GEN_960; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_962 = 10'h3c2 == csr_addr[9:0] ? reg_csr_962 : _GEN_961; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_963 = 10'h3c3 == csr_addr[9:0] ? reg_csr_963 : _GEN_962; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_964 = 10'h3c4 == csr_addr[9:0] ? reg_csr_964 : _GEN_963; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_965 = 10'h3c5 == csr_addr[9:0] ? reg_csr_965 : _GEN_964; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_966 = 10'h3c6 == csr_addr[9:0] ? reg_csr_966 : _GEN_965; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_967 = 10'h3c7 == csr_addr[9:0] ? reg_csr_967 : _GEN_966; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_968 = 10'h3c8 == csr_addr[9:0] ? reg_csr_968 : _GEN_967; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_969 = 10'h3c9 == csr_addr[9:0] ? reg_csr_969 : _GEN_968; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_970 = 10'h3ca == csr_addr[9:0] ? reg_csr_970 : _GEN_969; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_971 = 10'h3cb == csr_addr[9:0] ? reg_csr_971 : _GEN_970; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_972 = 10'h3cc == csr_addr[9:0] ? reg_csr_972 : _GEN_971; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_973 = 10'h3cd == csr_addr[9:0] ? reg_csr_973 : _GEN_972; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_974 = 10'h3ce == csr_addr[9:0] ? reg_csr_974 : _GEN_973; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_975 = 10'h3cf == csr_addr[9:0] ? reg_csr_975 : _GEN_974; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_976 = 10'h3d0 == csr_addr[9:0] ? reg_csr_976 : _GEN_975; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_977 = 10'h3d1 == csr_addr[9:0] ? reg_csr_977 : _GEN_976; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_978 = 10'h3d2 == csr_addr[9:0] ? reg_csr_978 : _GEN_977; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_979 = 10'h3d3 == csr_addr[9:0] ? reg_csr_979 : _GEN_978; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_980 = 10'h3d4 == csr_addr[9:0] ? reg_csr_980 : _GEN_979; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_981 = 10'h3d5 == csr_addr[9:0] ? reg_csr_981 : _GEN_980; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_982 = 10'h3d6 == csr_addr[9:0] ? reg_csr_982 : _GEN_981; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_983 = 10'h3d7 == csr_addr[9:0] ? reg_csr_983 : _GEN_982; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_984 = 10'h3d8 == csr_addr[9:0] ? reg_csr_984 : _GEN_983; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_985 = 10'h3d9 == csr_addr[9:0] ? reg_csr_985 : _GEN_984; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_986 = 10'h3da == csr_addr[9:0] ? reg_csr_986 : _GEN_985; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_987 = 10'h3db == csr_addr[9:0] ? reg_csr_987 : _GEN_986; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_988 = 10'h3dc == csr_addr[9:0] ? reg_csr_988 : _GEN_987; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_989 = 10'h3dd == csr_addr[9:0] ? reg_csr_989 : _GEN_988; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_990 = 10'h3de == csr_addr[9:0] ? reg_csr_990 : _GEN_989; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_991 = 10'h3df == csr_addr[9:0] ? reg_csr_991 : _GEN_990; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_992 = 10'h3e0 == csr_addr[9:0] ? reg_csr_992 : _GEN_991; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_993 = 10'h3e1 == csr_addr[9:0] ? reg_csr_993 : _GEN_992; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_994 = 10'h3e2 == csr_addr[9:0] ? reg_csr_994 : _GEN_993; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_995 = 10'h3e3 == csr_addr[9:0] ? reg_csr_995 : _GEN_994; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_996 = 10'h3e4 == csr_addr[9:0] ? reg_csr_996 : _GEN_995; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_997 = 10'h3e5 == csr_addr[9:0] ? reg_csr_997 : _GEN_996; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_998 = 10'h3e6 == csr_addr[9:0] ? reg_csr_998 : _GEN_997; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_999 = 10'h3e7 == csr_addr[9:0] ? reg_csr_999 : _GEN_998; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1000 = 10'h3e8 == csr_addr[9:0] ? reg_csr_1000 : _GEN_999; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1001 = 10'h3e9 == csr_addr[9:0] ? reg_csr_1001 : _GEN_1000; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1002 = 10'h3ea == csr_addr[9:0] ? reg_csr_1002 : _GEN_1001; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1003 = 10'h3eb == csr_addr[9:0] ? reg_csr_1003 : _GEN_1002; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1004 = 10'h3ec == csr_addr[9:0] ? reg_csr_1004 : _GEN_1003; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1005 = 10'h3ed == csr_addr[9:0] ? reg_csr_1005 : _GEN_1004; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1006 = 10'h3ee == csr_addr[9:0] ? reg_csr_1006 : _GEN_1005; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1007 = 10'h3ef == csr_addr[9:0] ? reg_csr_1007 : _GEN_1006; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1008 = 10'h3f0 == csr_addr[9:0] ? reg_csr_1008 : _GEN_1007; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1009 = 10'h3f1 == csr_addr[9:0] ? reg_csr_1009 : _GEN_1008; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1010 = 10'h3f2 == csr_addr[9:0] ? reg_csr_1010 : _GEN_1009; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1011 = 10'h3f3 == csr_addr[9:0] ? reg_csr_1011 : _GEN_1010; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1012 = 10'h3f4 == csr_addr[9:0] ? reg_csr_1012 : _GEN_1011; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1013 = 10'h3f5 == csr_addr[9:0] ? reg_csr_1013 : _GEN_1012; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1014 = 10'h3f6 == csr_addr[9:0] ? reg_csr_1014 : _GEN_1013; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1015 = 10'h3f7 == csr_addr[9:0] ? reg_csr_1015 : _GEN_1014; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1016 = 10'h3f8 == csr_addr[9:0] ? reg_csr_1016 : _GEN_1015; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1017 = 10'h3f9 == csr_addr[9:0] ? reg_csr_1017 : _GEN_1016; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1018 = 10'h3fa == csr_addr[9:0] ? reg_csr_1018 : _GEN_1017; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1019 = 10'h3fb == csr_addr[9:0] ? reg_csr_1019 : _GEN_1018; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1020 = 10'h3fc == csr_addr[9:0] ? reg_csr_1020 : _GEN_1019; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1021 = 10'h3fd == csr_addr[9:0] ? reg_csr_1021 : _GEN_1020; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1022 = 10'h3fe == csr_addr[9:0] ? reg_csr_1022 : _GEN_1021; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _GEN_1023 = 10'h3ff == csr_addr[9:0] ? reg_csr_1023 : _GEN_1022; // @[MEM.scala 83:43 MEM.scala 83:43]
  wire [31:0] _csr_wdata_T_2 = _GEN_1023 | io_in_id_in_op1_data; // @[MEM.scala 83:43]
  wire  _csr_wdata_T_3 = io_in_id_in_csr_cmd == 3'h3; // @[MEM.scala 84:18]
  wire [31:0] _csr_wdata_T_4 = ~io_in_id_in_op1_data; // @[MEM.scala 84:45]
  wire [31:0] _csr_wdata_T_5 = _GEN_1023 & _csr_wdata_T_4; // @[MEM.scala 84:43]
  wire [31:0] _csr_wdata_T_7 = _csr_addr_T ? 32'hb : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _csr_wdata_T_8 = _csr_wdata_T_3 ? _csr_wdata_T_5 : _csr_wdata_T_7; // @[Mux.scala 98:16]
  wire [31:0] _csr_wdata_T_9 = _csr_wdata_T_1 ? _csr_wdata_T_2 : _csr_wdata_T_8; // @[Mux.scala 98:16]
  wire [31:0] csr_wdata = _csr_wdata_T ? io_in_id_in_op1_data : _csr_wdata_T_9; // @[Mux.scala 98:16]
  wire  _rd_data_T = io_in_id_in_rd_sel == 3'h1; // @[MEM.scala 93:17]
  wire  _rd_data_T_1 = io_in_id_in_rd_sel == 3'h2; // @[MEM.scala 94:17]
  wire [31:0] _rd_data_T_3 = io_in_if_in_reg_pc + 32'h4; // @[MEM.scala 94:40]
  wire  _rd_data_T_4 = io_in_id_in_rd_sel == 3'h3; // @[MEM.scala 95:17]
  wire [31:0] _rd_data_T_5 = _rd_data_T_4 ? _GEN_1023 : io_in_ex_in_alu_out; // @[Mux.scala 98:16]
  wire [31:0] _rd_data_T_6 = _rd_data_T_1 ? _rd_data_T_3 : _rd_data_T_5; // @[Mux.scala 98:16]
  wire  _T_3 = ~reset; // @[MEM.scala 106:11]
  assign io_out_rd_wen = io_in_id_in_rd_wen; // @[MEM.scala 101:21]
  assign io_out_rd_addr = io_in_id_in_rd_addr; // @[MEM.scala 102:21]
  assign io_out_rd_data = _rd_data_T ? io_datamem_rdata : _rd_data_T_6; // @[Mux.scala 98:16]
  assign io_datamem_addr = io_in_ex_in_alu_out; // @[MEM.scala 72:25]
  assign io_datamem_wen = io_in_id_in_mem_wen; // @[MEM.scala 73:42]
  assign io_datamem_wdata = io_in_id_in_rs2_data; // @[MEM.scala 74:25]
  always @(posedge clock) begin
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_0 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_0 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_0 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_2 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_2 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_3 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_3 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_4 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_4 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_5 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_5 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_5 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_6 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_6 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_6 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_7 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_7 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_7 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_8 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_8 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_8 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_9 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_9 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_9 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_10 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_10 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_10 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_11 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_11 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_11 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_12 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_12 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_12 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_13 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_13 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_13 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_14 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_14 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_14 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_15 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_15 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_15 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_16 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_16 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_16 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_17 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_17 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_17 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_18 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_18 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_18 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_19 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_19 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_19 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_20 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_20 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_20 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_21 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_21 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_21 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_22 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_22 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_22 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_23 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_23 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_23 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_24 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_24 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_24 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_25 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_25 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_25 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_26 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_26 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_26 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_27 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_27 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_27 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_28 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_28 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_28 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_29 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_29 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_29 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_30 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_30 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_30 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_31 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_31 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_31 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_32 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_32 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_32 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_33 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_33 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_33 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_34 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_34 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_34 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_35 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_35 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_35 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_36 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_36 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_36 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_37 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_37 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_37 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_38 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_38 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_38 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_39 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_39 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_39 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_40 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_40 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_40 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_41 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_41 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_41 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_42 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_42 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_42 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_43 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_43 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_43 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_44 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_44 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_44 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_45 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_45 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_45 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_46 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_46 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_46 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_47 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_47 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_47 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_48 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_48 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_48 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_49 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_49 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_49 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_50 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_50 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_50 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_51 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_51 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_51 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_52 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_52 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_52 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_53 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_53 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_53 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_54 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_54 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_54 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_55 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_55 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_55 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_56 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_56 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_56 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_57 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_57 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_57 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_58 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_58 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_58 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_59 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_59 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_59 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_60 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_60 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_60 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_61 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_61 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_61 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_62 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_62 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_62 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_63 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_63 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_63 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_64 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h40 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_64 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_64 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_65 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h41 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_65 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_65 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_66 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h42 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_66 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_66 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_67 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h43 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_67 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_67 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_68 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h44 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_68 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_68 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_69 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h45 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_69 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_69 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_70 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h46 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_70 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_70 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_71 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h47 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_71 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_71 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_72 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h48 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_72 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_72 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_73 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h49 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_73 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_73 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_74 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_74 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_74 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_75 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_75 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_75 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_76 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_76 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_76 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_77 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_77 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_77 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_78 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_78 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_78 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_79 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h4f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_79 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_79 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_80 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h50 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_80 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_80 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_81 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h51 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_81 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_81 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_82 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h52 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_82 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_82 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_83 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h53 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_83 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_83 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_84 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h54 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_84 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_84 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_85 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h55 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_85 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_85 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_86 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h56 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_86 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_86 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_87 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h57 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_87 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_87 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_88 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h58 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_88 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_88 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_89 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h59 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_89 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_89 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_90 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_90 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_90 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_91 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_91 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_91 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_92 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_92 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_92 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_93 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_93 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_93 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_94 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_94 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_94 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_95 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h5f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_95 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_95 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_96 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h60 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_96 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_96 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_97 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h61 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_97 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_97 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_98 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h62 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_98 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_98 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_99 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h63 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_99 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_99 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_100 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h64 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_100 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_100 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_101 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h65 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_101 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_101 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_102 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h66 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_102 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_102 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_103 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h67 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_103 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_103 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_104 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h68 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_104 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_104 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_105 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h69 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_105 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_105 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_106 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_106 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_106 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_107 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_107 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_107 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_108 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_108 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_108 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_109 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_109 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_109 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_110 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_110 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_110 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_111 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h6f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_111 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_111 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_112 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h70 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_112 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_112 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_113 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h71 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_113 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_113 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_114 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h72 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_114 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_114 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_115 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h73 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_115 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_115 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_116 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h74 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_116 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_116 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_117 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h75 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_117 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_117 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_118 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h76 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_118 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_118 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_119 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h77 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_119 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_119 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_120 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h78 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_120 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_120 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_121 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h79 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_121 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_121 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_122 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_122 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_122 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_123 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_123 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_123 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_124 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_124 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_124 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_125 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_125 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_125 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_126 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_126 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_126 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_127 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h7f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_127 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_127 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_128 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h80 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_128 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_128 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_129 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h81 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_129 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_129 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_130 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h82 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_130 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_130 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_131 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h83 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_131 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_131 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_132 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h84 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_132 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_132 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_133 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h85 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_133 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_133 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_134 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h86 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_134 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_134 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_135 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h87 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_135 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_135 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_136 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h88 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_136 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_136 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_137 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h89 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_137 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_137 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_138 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_138 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_138 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_139 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_139 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_139 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_140 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_140 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_140 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_141 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_141 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_141 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_142 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_142 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_142 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_143 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h8f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_143 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_143 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_144 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h90 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_144 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_144 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_145 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h91 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_145 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_145 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_146 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h92 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_146 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_146 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_147 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h93 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_147 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_147 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_148 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h94 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_148 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_148 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_149 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h95 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_149 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_149 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_150 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h96 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_150 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_150 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_151 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h97 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_151 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_151 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_152 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h98 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_152 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_152 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_153 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h99 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_153 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_153 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_154 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_154 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_154 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_155 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_155 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_155 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_156 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_156 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_156 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_157 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_157 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_157 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_158 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_158 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_158 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_159 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h9f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_159 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_159 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_160 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_160 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_160 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_161 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_161 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_161 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_162 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_162 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_162 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_163 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_163 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_163 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_164 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_164 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_164 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_165 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_165 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_165 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_166 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_166 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_166 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_167 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_167 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_167 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_168 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_168 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_168 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_169 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'ha9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_169 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_169 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_170 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'haa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_170 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_170 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_171 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hab == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_171 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_171 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_172 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hac == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_172 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_172 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_173 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'had == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_173 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_173 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_174 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hae == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_174 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_174 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_175 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'haf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_175 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_175 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_176 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_176 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_176 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_177 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_177 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_177 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_178 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_178 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_178 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_179 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_179 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_179 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_180 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_180 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_180 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_181 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_181 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_181 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_182 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_182 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_182 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_183 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_183 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_183 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_184 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_184 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_184 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_185 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hb9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_185 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_185 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_186 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hba == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_186 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_186 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_187 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hbb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_187 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_187 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_188 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hbc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_188 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_188 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_189 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hbd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_189 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_189 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_190 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hbe == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_190 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_190 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_191 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hbf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_191 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_191 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_192 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_192 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_192 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_193 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_193 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_193 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_194 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_194 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_194 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_195 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_195 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_195 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_196 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_196 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_196 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_197 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_197 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_197 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_198 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_198 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_198 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_199 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_199 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_199 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_200 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_200 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_200 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_201 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hc9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_201 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_201 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_202 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hca == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_202 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_202 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_203 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hcb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_203 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_203 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_204 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hcc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_204 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_204 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_205 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hcd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_205 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_205 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_206 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hce == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_206 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_206 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_207 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hcf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_207 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_207 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_208 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_208 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_208 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_209 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_209 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_209 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_210 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_210 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_210 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_211 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_211 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_211 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_212 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_212 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_212 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_213 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_213 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_213 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_214 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_214 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_214 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_215 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_215 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_215 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_216 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_216 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_216 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_217 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hd9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_217 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_217 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_218 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hda == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_218 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_218 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_219 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hdb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_219 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_219 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_220 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hdc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_220 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_220 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_221 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hdd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_221 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_221 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_222 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hde == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_222 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_222 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_223 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hdf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_223 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_223 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_224 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_224 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_224 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_225 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_225 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_225 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_226 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_226 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_226 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_227 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_227 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_227 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_228 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_228 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_228 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_229 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_229 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_229 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_230 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_230 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_230 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_231 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_231 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_231 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_232 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_232 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_232 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_233 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'he9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_233 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_233 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_234 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hea == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_234 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_234 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_235 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'heb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_235 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_235 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_236 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hec == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_236 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_236 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_237 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hed == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_237 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_237 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_238 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hee == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_238 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_238 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_239 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hef == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_239 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_239 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_240 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_240 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_240 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_241 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_241 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_241 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_242 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_242 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_242 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_243 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_243 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_243 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_244 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_244 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_244 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_245 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_245 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_245 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_246 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_246 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_246 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_247 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_247 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_247 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_248 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_248 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_248 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_249 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hf9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_249 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_249 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_250 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hfa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_250 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_250 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_251 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hfb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_251 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_251 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_252 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hfc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_252 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_252 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_253 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hfd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_253 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_253 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_254 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hfe == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_254 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_254 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_255 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'hff == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_255 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_255 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_256 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h100 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_256 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_256 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_257 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h101 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_257 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_257 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_258 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h102 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_258 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_258 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_259 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h103 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_259 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_259 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_260 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h104 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_260 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_260 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_261 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h105 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_261 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_261 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_262 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h106 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_262 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_262 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_263 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h107 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_263 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_263 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_264 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h108 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_264 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_264 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_265 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h109 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_265 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_265 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_266 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_266 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_266 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_267 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_267 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_267 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_268 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_268 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_268 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_269 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_269 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_269 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_270 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_270 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_270 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_271 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h10f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_271 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_271 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_272 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h110 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_272 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_272 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_273 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h111 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_273 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_273 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_274 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h112 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_274 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_274 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_275 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h113 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_275 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_275 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_276 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h114 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_276 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_276 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_277 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h115 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_277 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_277 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_278 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h116 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_278 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_278 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_279 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h117 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_279 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_279 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_280 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h118 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_280 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_280 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_281 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h119 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_281 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_281 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_282 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_282 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_282 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_283 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_283 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_283 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_284 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_284 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_284 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_285 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_285 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_285 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_286 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_286 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_286 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_287 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h11f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_287 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_287 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_288 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h120 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_288 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_288 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_289 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h121 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_289 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_289 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_290 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h122 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_290 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_290 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_291 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h123 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_291 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_291 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_292 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h124 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_292 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_292 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_293 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h125 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_293 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_293 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_294 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h126 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_294 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_294 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_295 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h127 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_295 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_295 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_296 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h128 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_296 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_296 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_297 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h129 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_297 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_297 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_298 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_298 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_298 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_299 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_299 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_299 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_300 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_300 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_300 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_301 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_301 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_301 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_302 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_302 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_302 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_303 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h12f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_303 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_303 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_304 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h130 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_304 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_304 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_305 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h131 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_305 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_305 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_306 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h132 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_306 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_306 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_307 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h133 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_307 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_307 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_308 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h134 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_308 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_308 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_309 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h135 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_309 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_309 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_310 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h136 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_310 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_310 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_311 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h137 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_311 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_311 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_312 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h138 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_312 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_312 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_313 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h139 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_313 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_313 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_314 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_314 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_314 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_315 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_315 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_315 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_316 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_316 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_316 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_317 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_317 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_317 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_318 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_318 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_318 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_319 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h13f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_319 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_319 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_320 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h140 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_320 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_320 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_321 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h141 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_321 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_321 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_322 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h142 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_322 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_322 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_323 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h143 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_323 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_323 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_324 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h144 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_324 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_324 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_325 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h145 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_325 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_325 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_326 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h146 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_326 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_326 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_327 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h147 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_327 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_327 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_328 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h148 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_328 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_328 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_329 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h149 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_329 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_329 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_330 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_330 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_330 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_331 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_331 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_331 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_332 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_332 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_332 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_333 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_333 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_333 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_334 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_334 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_334 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_335 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h14f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_335 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_335 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_336 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h150 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_336 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_336 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_337 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h151 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_337 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_337 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_338 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h152 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_338 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_338 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_339 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h153 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_339 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_339 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_340 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h154 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_340 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_340 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_341 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h155 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_341 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_341 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_342 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h156 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_342 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_342 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_343 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h157 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_343 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_343 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_344 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h158 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_344 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_344 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_345 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h159 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_345 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_345 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_346 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_346 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_346 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_347 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_347 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_347 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_348 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_348 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_348 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_349 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_349 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_349 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_350 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_350 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_350 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_351 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h15f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_351 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_351 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_352 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h160 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_352 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_352 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_353 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h161 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_353 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_353 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_354 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h162 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_354 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_354 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_355 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h163 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_355 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_355 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_356 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h164 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_356 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_356 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_357 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h165 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_357 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_357 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_358 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h166 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_358 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_358 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_359 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h167 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_359 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_359 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_360 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h168 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_360 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_360 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_361 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h169 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_361 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_361 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_362 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_362 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_362 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_363 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_363 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_363 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_364 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_364 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_364 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_365 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_365 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_365 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_366 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_366 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_366 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_367 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h16f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_367 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_367 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_368 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h170 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_368 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_368 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_369 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h171 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_369 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_369 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_370 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h172 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_370 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_370 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_371 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h173 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_371 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_371 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_372 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h174 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_372 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_372 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_373 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h175 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_373 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_373 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_374 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h176 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_374 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_374 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_375 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h177 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_375 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_375 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_376 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h178 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_376 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_376 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_377 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h179 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_377 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_377 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_378 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_378 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_378 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_379 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_379 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_379 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_380 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_380 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_380 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_381 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_381 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_381 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_382 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_382 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_382 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_383 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h17f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_383 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_383 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_384 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h180 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_384 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_384 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_385 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h181 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_385 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_385 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_386 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h182 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_386 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_386 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_387 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h183 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_387 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_387 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_388 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h184 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_388 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_388 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_389 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h185 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_389 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_389 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_390 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h186 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_390 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_390 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_391 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h187 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_391 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_391 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_392 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h188 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_392 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_392 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_393 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h189 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_393 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_393 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_394 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_394 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_394 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_395 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_395 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_395 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_396 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_396 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_396 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_397 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_397 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_397 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_398 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_398 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_398 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_399 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h18f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_399 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_399 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_400 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h190 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_400 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_400 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_401 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h191 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_401 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_401 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_402 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h192 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_402 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_402 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_403 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h193 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_403 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_403 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_404 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h194 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_404 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_404 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_405 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h195 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_405 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_405 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_406 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h196 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_406 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_406 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_407 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h197 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_407 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_407 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_408 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h198 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_408 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_408 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_409 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h199 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_409 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_409 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_410 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_410 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_410 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_411 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_411 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_411 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_412 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_412 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_412 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_413 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_413 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_413 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_414 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_414 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_414 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_415 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h19f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_415 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_415 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_416 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_416 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_416 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_417 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_417 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_417 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_418 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_418 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_418 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_419 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_419 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_419 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_420 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_420 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_420 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_421 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_421 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_421 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_422 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_422 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_422 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_423 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_423 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_423 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_424 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_424 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_424 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_425 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1a9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_425 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_425 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_426 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1aa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_426 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_426 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_427 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ab == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_427 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_427 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_428 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ac == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_428 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_428 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_429 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ad == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_429 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_429 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_430 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ae == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_430 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_430 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_431 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1af == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_431 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_431 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_432 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_432 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_432 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_433 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_433 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_433 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_434 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_434 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_434 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_435 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_435 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_435 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_436 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_436 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_436 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_437 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_437 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_437 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_438 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_438 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_438 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_439 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_439 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_439 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_440 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_440 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_440 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_441 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1b9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_441 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_441 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_442 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ba == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_442 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_442 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_443 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1bb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_443 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_443 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_444 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1bc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_444 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_444 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_445 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1bd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_445 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_445 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_446 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1be == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_446 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_446 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_447 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1bf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_447 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_447 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_448 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_448 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_448 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_449 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_449 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_449 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_450 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_450 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_450 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_451 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_451 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_451 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_452 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_452 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_452 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_453 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_453 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_453 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_454 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_454 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_454 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_455 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_455 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_455 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_456 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_456 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_456 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_457 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1c9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_457 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_457 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_458 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ca == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_458 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_458 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_459 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1cb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_459 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_459 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_460 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1cc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_460 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_460 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_461 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1cd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_461 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_461 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_462 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ce == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_462 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_462 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_463 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1cf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_463 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_463 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_464 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_464 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_464 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_465 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_465 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_465 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_466 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_466 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_466 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_467 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_467 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_467 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_468 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_468 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_468 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_469 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_469 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_469 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_470 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_470 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_470 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_471 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_471 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_471 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_472 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_472 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_472 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_473 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1d9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_473 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_473 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_474 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1da == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_474 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_474 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_475 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1db == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_475 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_475 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_476 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1dc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_476 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_476 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_477 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1dd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_477 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_477 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_478 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1de == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_478 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_478 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_479 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1df == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_479 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_479 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_480 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_480 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_480 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_481 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_481 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_481 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_482 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_482 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_482 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_483 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_483 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_483 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_484 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_484 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_484 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_485 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_485 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_485 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_486 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_486 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_486 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_487 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_487 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_487 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_488 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_488 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_488 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_489 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1e9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_489 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_489 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_490 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ea == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_490 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_490 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_491 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1eb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_491 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_491 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_492 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ec == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_492 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_492 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_493 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ed == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_493 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_493 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_494 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ee == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_494 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_494 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_495 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ef == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_495 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_495 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_496 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_496 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_496 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_497 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_497 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_497 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_498 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_498 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_498 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_499 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_499 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_499 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_500 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_500 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_500 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_501 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_501 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_501 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_502 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_502 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_502 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_503 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_503 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_503 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_504 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_504 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_504 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_505 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1f9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_505 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_505 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_506 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1fa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_506 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_506 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_507 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1fb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_507 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_507 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_508 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1fc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_508 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_508 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_509 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1fd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_509 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_509 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_510 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1fe == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_510 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_510 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_511 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h1ff == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_511 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_511 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_512 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h200 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_512 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_512 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_513 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h201 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_513 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_513 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_514 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h202 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_514 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_514 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_515 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h203 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_515 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_515 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_516 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h204 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_516 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_516 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_517 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h205 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_517 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_517 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_518 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h206 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_518 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_518 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_519 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h207 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_519 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_519 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_520 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h208 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_520 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_520 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_521 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h209 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_521 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_521 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_522 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_522 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_522 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_523 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_523 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_523 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_524 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_524 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_524 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_525 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_525 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_525 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_526 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_526 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_526 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_527 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h20f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_527 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_527 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_528 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h210 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_528 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_528 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_529 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h211 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_529 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_529 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_530 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h212 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_530 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_530 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_531 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h213 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_531 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_531 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_532 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h214 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_532 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_532 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_533 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h215 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_533 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_533 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_534 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h216 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_534 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_534 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_535 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h217 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_535 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_535 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_536 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h218 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_536 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_536 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_537 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h219 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_537 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_537 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_538 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_538 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_538 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_539 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_539 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_539 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_540 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_540 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_540 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_541 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_541 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_541 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_542 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_542 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_542 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_543 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h21f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_543 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_543 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_544 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h220 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_544 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_544 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_545 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h221 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_545 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_545 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_546 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h222 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_546 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_546 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_547 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h223 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_547 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_547 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_548 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h224 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_548 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_548 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_549 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h225 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_549 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_549 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_550 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h226 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_550 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_550 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_551 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h227 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_551 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_551 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_552 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h228 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_552 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_552 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_553 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h229 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_553 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_553 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_554 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_554 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_554 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_555 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_555 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_555 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_556 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_556 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_556 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_557 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_557 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_557 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_558 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_558 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_558 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_559 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h22f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_559 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_559 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_560 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h230 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_560 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_560 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_561 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h231 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_561 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_561 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_562 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h232 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_562 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_562 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_563 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h233 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_563 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_563 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_564 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h234 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_564 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_564 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_565 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h235 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_565 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_565 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_566 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h236 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_566 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_566 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_567 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h237 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_567 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_567 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_568 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h238 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_568 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_568 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_569 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h239 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_569 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_569 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_570 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_570 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_570 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_571 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_571 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_571 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_572 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_572 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_572 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_573 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_573 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_573 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_574 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_574 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_574 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_575 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h23f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_575 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_575 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_576 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h240 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_576 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_576 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_577 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h241 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_577 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_577 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_578 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h242 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_578 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_578 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_579 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h243 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_579 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_579 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_580 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h244 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_580 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_580 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_581 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h245 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_581 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_581 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_582 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h246 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_582 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_582 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_583 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h247 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_583 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_583 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_584 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h248 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_584 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_584 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_585 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h249 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_585 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_585 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_586 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_586 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_586 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_587 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_587 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_587 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_588 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_588 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_588 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_589 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_589 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_589 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_590 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_590 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_590 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_591 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h24f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_591 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_591 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_592 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h250 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_592 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_592 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_593 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h251 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_593 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_593 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_594 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h252 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_594 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_594 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_595 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h253 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_595 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_595 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_596 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h254 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_596 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_596 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_597 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h255 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_597 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_597 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_598 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h256 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_598 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_598 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_599 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h257 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_599 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_599 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_600 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h258 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_600 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_600 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_601 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h259 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_601 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_601 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_602 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_602 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_602 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_603 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_603 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_603 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_604 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_604 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_604 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_605 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_605 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_605 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_606 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_606 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_606 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_607 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h25f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_607 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_607 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_608 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h260 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_608 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_608 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_609 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h261 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_609 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_609 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_610 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h262 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_610 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_610 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_611 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h263 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_611 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_611 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_612 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h264 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_612 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_612 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_613 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h265 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_613 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_613 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_614 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h266 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_614 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_614 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_615 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h267 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_615 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_615 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_616 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h268 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_616 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_616 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_617 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h269 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_617 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_617 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_618 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_618 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_618 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_619 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_619 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_619 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_620 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_620 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_620 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_621 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_621 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_621 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_622 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_622 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_622 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_623 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h26f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_623 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_623 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_624 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h270 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_624 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_624 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_625 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h271 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_625 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_625 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_626 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h272 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_626 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_626 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_627 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h273 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_627 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_627 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_628 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h274 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_628 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_628 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_629 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h275 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_629 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_629 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_630 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h276 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_630 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_630 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_631 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h277 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_631 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_631 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_632 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h278 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_632 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_632 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_633 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h279 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_633 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_633 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_634 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_634 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_634 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_635 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_635 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_635 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_636 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_636 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_636 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_637 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_637 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_637 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_638 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_638 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_638 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_639 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h27f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_639 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_639 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_640 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h280 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_640 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_640 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_641 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h281 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_641 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_641 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_642 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h282 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_642 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_642 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_643 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h283 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_643 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_643 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_644 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h284 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_644 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_644 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_645 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h285 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_645 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_645 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_646 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h286 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_646 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_646 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_647 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h287 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_647 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_647 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_648 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h288 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_648 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_648 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_649 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h289 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_649 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_649 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_650 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_650 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_650 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_651 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_651 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_651 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_652 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_652 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_652 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_653 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_653 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_653 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_654 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_654 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_654 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_655 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h28f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_655 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_655 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_656 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h290 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_656 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_656 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_657 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h291 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_657 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_657 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_658 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h292 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_658 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_658 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_659 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h293 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_659 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_659 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_660 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h294 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_660 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_660 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_661 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h295 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_661 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_661 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_662 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h296 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_662 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_662 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_663 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h297 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_663 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_663 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_664 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h298 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_664 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_664 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_665 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h299 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_665 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_665 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_666 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_666 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_666 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_667 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_667 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_667 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_668 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_668 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_668 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_669 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_669 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_669 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_670 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_670 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_670 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_671 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h29f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_671 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_671 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_672 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_672 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_672 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_673 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_673 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_673 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_674 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_674 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_674 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_675 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_675 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_675 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_676 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_676 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_676 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_677 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_677 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_677 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_678 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_678 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_678 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_679 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_679 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_679 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_680 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_680 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_680 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_681 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2a9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_681 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_681 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_682 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2aa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_682 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_682 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_683 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ab == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_683 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_683 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_684 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ac == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_684 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_684 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_685 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ad == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_685 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_685 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_686 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ae == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_686 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_686 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_687 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2af == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_687 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_687 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_688 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_688 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_688 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_689 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_689 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_689 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_690 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_690 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_690 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_691 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_691 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_691 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_692 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_692 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_692 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_693 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_693 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_693 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_694 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_694 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_694 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_695 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_695 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_695 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_696 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_696 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_696 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_697 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2b9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_697 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_697 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_698 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ba == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_698 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_698 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_699 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2bb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_699 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_699 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_700 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2bc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_700 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_700 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_701 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2bd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_701 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_701 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_702 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2be == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_702 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_702 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_703 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2bf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_703 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_703 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_704 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_704 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_704 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_705 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_705 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_705 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_706 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_706 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_706 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_707 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_707 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_707 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_708 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_708 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_708 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_709 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_709 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_709 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_710 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_710 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_710 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_711 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_711 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_711 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_712 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_712 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_712 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_713 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2c9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_713 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_713 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_714 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ca == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_714 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_714 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_715 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2cb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_715 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_715 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_716 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2cc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_716 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_716 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_717 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2cd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_717 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_717 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_718 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ce == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_718 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_718 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_719 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2cf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_719 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_719 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_720 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_720 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_720 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_721 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_721 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_721 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_722 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_722 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_722 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_723 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_723 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_723 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_724 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_724 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_724 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_725 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_725 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_725 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_726 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_726 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_726 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_727 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_727 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_727 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_728 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_728 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_728 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_729 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2d9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_729 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_729 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_730 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2da == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_730 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_730 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_731 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2db == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_731 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_731 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_732 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2dc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_732 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_732 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_733 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2dd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_733 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_733 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_734 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2de == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_734 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_734 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_735 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2df == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_735 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_735 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_736 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_736 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_736 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_737 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_737 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_737 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_738 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_738 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_738 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_739 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_739 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_739 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_740 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_740 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_740 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_741 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_741 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_741 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_742 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_742 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_742 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_743 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_743 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_743 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_744 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_744 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_744 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_745 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2e9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_745 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_745 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_746 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ea == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_746 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_746 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_747 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2eb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_747 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_747 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_748 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ec == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_748 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_748 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_749 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ed == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_749 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_749 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_750 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ee == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_750 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_750 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_751 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ef == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_751 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_751 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_752 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_752 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_752 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_753 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_753 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_753 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_754 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_754 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_754 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_755 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_755 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_755 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_756 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_756 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_756 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_757 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_757 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_757 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_758 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_758 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_758 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_759 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_759 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_759 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_760 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_760 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_760 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_761 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2f9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_761 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_761 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_762 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2fa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_762 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_762 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_763 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2fb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_763 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_763 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_764 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2fc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_764 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_764 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_765 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2fd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_765 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_765 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_766 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2fe == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_766 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_766 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_767 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h2ff == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_767 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_767 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_768 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h300 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_768 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_768 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_769 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h301 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_769 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_769 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_770 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h302 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_770 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_770 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_771 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h303 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_771 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_771 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_772 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h304 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_772 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_772 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_773 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h305 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_773 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_773 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_774 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h306 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_774 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_774 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_775 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h307 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_775 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_775 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_776 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h308 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_776 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_776 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_777 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h309 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_777 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_777 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_778 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_778 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_778 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_779 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_779 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_779 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_780 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_780 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_780 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_781 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_781 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_781 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_782 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_782 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_782 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_783 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h30f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_783 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_783 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_784 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h310 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_784 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_784 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_785 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h311 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_785 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_785 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_786 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h312 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_786 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_786 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_787 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h313 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_787 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_787 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_788 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h314 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_788 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_788 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_789 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h315 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_789 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_789 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_790 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h316 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_790 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_790 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_791 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h317 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_791 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_791 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_792 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h318 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_792 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_792 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_793 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h319 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_793 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_793 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_794 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_794 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_794 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_795 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_795 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_795 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_796 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_796 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_796 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_797 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_797 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_797 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_798 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_798 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_798 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_799 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h31f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_799 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_799 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_800 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h320 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_800 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_800 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_801 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h321 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_801 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_801 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_802 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h322 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_802 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_802 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_803 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h323 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_803 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_803 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_804 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h324 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_804 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_804 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_805 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h325 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_805 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_805 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_806 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h326 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_806 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_806 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_807 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h327 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_807 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_807 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_808 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h328 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_808 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_808 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_809 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h329 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_809 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_809 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_810 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_810 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_810 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_811 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_811 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_811 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_812 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_812 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_812 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_813 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_813 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_813 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_814 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_814 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_814 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_815 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h32f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_815 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_815 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_816 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h330 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_816 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_816 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_817 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h331 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_817 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_817 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_818 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h332 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_818 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_818 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_819 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h333 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_819 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_819 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_820 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h334 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_820 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_820 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_821 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h335 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_821 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_821 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_822 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h336 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_822 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_822 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_823 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h337 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_823 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_823 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_824 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h338 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_824 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_824 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_825 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h339 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_825 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_825 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_826 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_826 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_826 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_827 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_827 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_827 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_828 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_828 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_828 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_829 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_829 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_829 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_830 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_830 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_830 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_831 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h33f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_831 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_831 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_832 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h340 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_832 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_832 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_833 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h341 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_833 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_833 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_834 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h342 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_834 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_834 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_835 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h343 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_835 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_835 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_836 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h344 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_836 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_836 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_837 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h345 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_837 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_837 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_838 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h346 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_838 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_838 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_839 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h347 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_839 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_839 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_840 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h348 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_840 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_840 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_841 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h349 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_841 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_841 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_842 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_842 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_842 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_843 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_843 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_843 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_844 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_844 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_844 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_845 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_845 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_845 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_846 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_846 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_846 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_847 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h34f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_847 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_847 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_848 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h350 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_848 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_848 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_849 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h351 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_849 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_849 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_850 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h352 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_850 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_850 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_851 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h353 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_851 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_851 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_852 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h354 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_852 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_852 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_853 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h355 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_853 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_853 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_854 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h356 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_854 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_854 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_855 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h357 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_855 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_855 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_856 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h358 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_856 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_856 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_857 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h359 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_857 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_857 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_858 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_858 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_858 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_859 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_859 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_859 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_860 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_860 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_860 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_861 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_861 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_861 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_862 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_862 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_862 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_863 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h35f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_863 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_863 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_864 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h360 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_864 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_864 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_865 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h361 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_865 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_865 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_866 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h362 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_866 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_866 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_867 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h363 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_867 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_867 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_868 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h364 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_868 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_868 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_869 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h365 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_869 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_869 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_870 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h366 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_870 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_870 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_871 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h367 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_871 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_871 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_872 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h368 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_872 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_872 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_873 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h369 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_873 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_873 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_874 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_874 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_874 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_875 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_875 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_875 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_876 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_876 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_876 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_877 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_877 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_877 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_878 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_878 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_878 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_879 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h36f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_879 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_879 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_880 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h370 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_880 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_880 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_881 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h371 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_881 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_881 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_882 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h372 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_882 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_882 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_883 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h373 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_883 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_883 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_884 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h374 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_884 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_884 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_885 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h375 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_885 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_885 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_886 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h376 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_886 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_886 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_887 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h377 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_887 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_887 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_888 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h378 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_888 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_888 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_889 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h379 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_889 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_889 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_890 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_890 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_890 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_891 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_891 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_891 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_892 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_892 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_892 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_893 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_893 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_893 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_894 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_894 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_894 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_895 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h37f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_895 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_895 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_896 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h380 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_896 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_896 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_897 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h381 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_897 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_897 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_898 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h382 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_898 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_898 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_899 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h383 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_899 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_899 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_900 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h384 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_900 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_900 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_901 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h385 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_901 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_901 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_902 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h386 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_902 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_902 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_903 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h387 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_903 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_903 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_904 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h388 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_904 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_904 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_905 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h389 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_905 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_905 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_906 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_906 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_906 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_907 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_907 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_907 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_908 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_908 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_908 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_909 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_909 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_909 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_910 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_910 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_910 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_911 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h38f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_911 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_911 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_912 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h390 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_912 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_912 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_913 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h391 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_913 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_913 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_914 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h392 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_914 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_914 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_915 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h393 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_915 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_915 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_916 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h394 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_916 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_916 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_917 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h395 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_917 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_917 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_918 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h396 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_918 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_918 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_919 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h397 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_919 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_919 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_920 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h398 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_920 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_920 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_921 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h399 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_921 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_921 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_922 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39a == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_922 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_922 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_923 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39b == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_923 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_923 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_924 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39c == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_924 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_924 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_925 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39d == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_925 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_925 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_926 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39e == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_926 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_926 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_927 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h39f == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_927 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_927 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_928 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_928 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_928 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_929 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_929 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_929 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_930 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_930 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_930 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_931 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_931 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_931 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_932 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_932 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_932 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_933 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_933 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_933 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_934 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_934 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_934 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_935 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_935 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_935 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_936 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_936 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_936 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_937 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3a9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_937 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_937 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_938 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3aa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_938 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_938 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_939 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ab == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_939 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_939 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_940 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ac == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_940 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_940 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_941 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ad == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_941 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_941 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_942 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ae == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_942 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_942 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_943 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3af == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_943 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_943 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_944 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_944 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_944 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_945 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_945 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_945 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_946 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_946 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_946 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_947 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_947 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_947 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_948 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_948 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_948 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_949 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_949 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_949 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_950 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_950 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_950 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_951 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_951 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_951 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_952 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_952 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_952 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_953 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3b9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_953 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_953 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_954 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ba == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_954 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_954 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_955 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3bb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_955 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_955 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_956 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3bc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_956 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_956 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_957 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3bd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_957 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_957 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_958 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3be == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_958 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_958 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_959 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3bf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_959 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_959 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_960 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_960 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_960 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_961 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_961 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_961 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_962 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_962 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_962 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_963 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_963 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_963 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_964 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_964 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_964 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_965 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_965 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_965 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_966 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_966 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_966 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_967 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_967 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_967 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_968 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_968 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_968 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_969 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3c9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_969 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_969 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_970 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ca == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_970 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_970 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_971 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3cb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_971 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_971 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_972 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3cc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_972 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_972 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_973 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3cd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_973 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_973 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_974 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ce == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_974 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_974 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_975 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3cf == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_975 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_975 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_976 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_976 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_976 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_977 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_977 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_977 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_978 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_978 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_978 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_979 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_979 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_979 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_980 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_980 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_980 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_981 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_981 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_981 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_982 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_982 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_982 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_983 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_983 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_983 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_984 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_984 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_984 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_985 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3d9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_985 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_985 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_986 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3da == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_986 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_986 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_987 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3db == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_987 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_987 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_988 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3dc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_988 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_988 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_989 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3dd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_989 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_989 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_990 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3de == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_990 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_990 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_991 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3df == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_991 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_991 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_992 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_992 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_992 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_993 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_993 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_993 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_994 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_994 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_994 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_995 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_995 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_995 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_996 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_996 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_996 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_997 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_997 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_997 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_998 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_998 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_998 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_999 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_999 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_999 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1000 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1000 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1000 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1001 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3e9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1001 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1001 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1002 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ea == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1002 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1002 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1003 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3eb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1003 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1003 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1004 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ec == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1004 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1004 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1005 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ed == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1005 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1005 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1006 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ee == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1006 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1006 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1007 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ef == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1007 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1007 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1008 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f0 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1008 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1008 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1009 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f1 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1009 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1009 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1010 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f2 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1010 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1010 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1011 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f3 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1011 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1011 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1012 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f4 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1012 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1012 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1013 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f5 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1013 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1013 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1014 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f6 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1014 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1014 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1015 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f7 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1015 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1015 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1016 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f8 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1016 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1016 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1017 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3f9 == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1017 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1017 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1018 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3fa == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1018 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1018 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1019 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3fb == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1019 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1019 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1020 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3fc == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1020 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1020 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1021 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3fd == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1021 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1021 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1022 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3fe == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1022 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1022 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[MEM.scala 54:26]
      reg_csr_1023 <= 32'h0; // @[MEM.scala 54:26]
    end else if (io_in_id_in_csr_cmd != 3'h0) begin // @[MEM.scala 87:31]
      if (10'h3ff == csr_addr[9:0]) begin // @[MEM.scala 88:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1023 <= io_in_id_in_op1_data;
        end else begin
          reg_csr_1023 <= _csr_wdata_T_9;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------MEM-----------\n"); // @[MEM.scala 106:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"datamem.wen: %d\n",io_datamem_wen); // @[MEM.scala 107:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"datamem.wdata: 0x%x\n",io_datamem_wdata); // @[MEM.scala 108:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"csr_wdata: 0x%x\n",csr_wdata); // @[MEM.scala 109:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_csr_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_csr_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_csr_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_csr_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_csr_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_csr_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_csr_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_csr_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_csr_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_csr_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_csr_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_csr_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_csr_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_csr_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_csr_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_csr_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_csr_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_csr_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_csr_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_csr_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_csr_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_csr_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_csr_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_csr_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_csr_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_csr_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_csr_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_csr_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_csr_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_csr_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_csr_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_csr_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  reg_csr_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  reg_csr_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  reg_csr_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  reg_csr_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_csr_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_csr_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_csr_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  reg_csr_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_csr_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  reg_csr_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  reg_csr_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  reg_csr_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  reg_csr_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  reg_csr_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  reg_csr_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  reg_csr_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_csr_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_csr_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  reg_csr_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  reg_csr_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  reg_csr_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  reg_csr_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  reg_csr_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  reg_csr_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  reg_csr_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  reg_csr_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  reg_csr_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  reg_csr_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  reg_csr_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  reg_csr_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  reg_csr_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  reg_csr_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  reg_csr_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  reg_csr_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  reg_csr_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  reg_csr_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  reg_csr_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  reg_csr_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  reg_csr_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  reg_csr_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  reg_csr_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  reg_csr_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  reg_csr_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  reg_csr_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  reg_csr_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  reg_csr_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  reg_csr_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  reg_csr_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  reg_csr_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  reg_csr_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  reg_csr_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  reg_csr_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  reg_csr_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  reg_csr_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  reg_csr_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  reg_csr_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  reg_csr_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  reg_csr_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  reg_csr_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  reg_csr_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  reg_csr_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  reg_csr_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  reg_csr_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  reg_csr_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  reg_csr_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  reg_csr_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  reg_csr_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  reg_csr_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  reg_csr_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  reg_csr_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  reg_csr_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  reg_csr_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  reg_csr_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  reg_csr_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  reg_csr_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  reg_csr_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  reg_csr_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  reg_csr_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  reg_csr_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  reg_csr_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  reg_csr_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  reg_csr_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  reg_csr_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  reg_csr_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  reg_csr_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  reg_csr_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  reg_csr_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  reg_csr_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  reg_csr_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  reg_csr_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  reg_csr_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  reg_csr_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  reg_csr_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  reg_csr_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  reg_csr_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  reg_csr_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  reg_csr_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  reg_csr_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  reg_csr_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  reg_csr_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  reg_csr_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  reg_csr_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  reg_csr_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  reg_csr_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  reg_csr_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  reg_csr_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  reg_csr_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  reg_csr_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  reg_csr_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  reg_csr_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  reg_csr_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  reg_csr_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  reg_csr_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  reg_csr_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  reg_csr_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  reg_csr_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  reg_csr_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  reg_csr_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  reg_csr_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  reg_csr_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  reg_csr_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  reg_csr_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  reg_csr_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  reg_csr_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  reg_csr_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  reg_csr_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  reg_csr_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  reg_csr_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  reg_csr_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  reg_csr_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  reg_csr_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  reg_csr_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  reg_csr_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  reg_csr_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  reg_csr_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  reg_csr_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  reg_csr_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  reg_csr_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  reg_csr_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  reg_csr_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  reg_csr_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  reg_csr_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  reg_csr_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  reg_csr_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  reg_csr_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  reg_csr_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  reg_csr_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  reg_csr_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  reg_csr_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  reg_csr_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  reg_csr_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  reg_csr_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  reg_csr_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  reg_csr_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  reg_csr_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  reg_csr_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  reg_csr_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  reg_csr_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  reg_csr_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  reg_csr_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  reg_csr_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  reg_csr_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  reg_csr_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  reg_csr_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  reg_csr_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  reg_csr_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  reg_csr_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  reg_csr_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  reg_csr_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  reg_csr_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  reg_csr_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  reg_csr_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  reg_csr_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  reg_csr_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  reg_csr_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  reg_csr_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  reg_csr_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  reg_csr_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  reg_csr_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  reg_csr_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  reg_csr_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  reg_csr_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  reg_csr_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  reg_csr_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  reg_csr_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  reg_csr_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  reg_csr_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  reg_csr_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  reg_csr_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  reg_csr_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  reg_csr_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  reg_csr_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  reg_csr_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  reg_csr_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  reg_csr_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  reg_csr_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  reg_csr_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  reg_csr_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  reg_csr_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  reg_csr_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  reg_csr_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  reg_csr_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  reg_csr_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  reg_csr_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  reg_csr_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  reg_csr_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  reg_csr_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  reg_csr_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  reg_csr_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  reg_csr_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  reg_csr_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  reg_csr_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  reg_csr_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  reg_csr_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  reg_csr_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  reg_csr_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  reg_csr_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  reg_csr_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  reg_csr_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  reg_csr_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  reg_csr_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  reg_csr_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  reg_csr_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  reg_csr_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  reg_csr_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  reg_csr_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  reg_csr_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  reg_csr_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  reg_csr_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  reg_csr_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  reg_csr_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  reg_csr_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  reg_csr_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  reg_csr_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  reg_csr_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  reg_csr_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  reg_csr_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  reg_csr_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  reg_csr_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  reg_csr_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  reg_csr_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  reg_csr_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  reg_csr_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  reg_csr_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  reg_csr_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  reg_csr_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  reg_csr_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  reg_csr_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  reg_csr_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  reg_csr_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  reg_csr_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  reg_csr_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  reg_csr_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  reg_csr_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  reg_csr_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  reg_csr_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  reg_csr_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  reg_csr_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  reg_csr_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  reg_csr_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  reg_csr_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  reg_csr_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  reg_csr_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  reg_csr_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  reg_csr_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  reg_csr_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  reg_csr_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  reg_csr_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  reg_csr_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  reg_csr_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  reg_csr_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  reg_csr_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  reg_csr_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  reg_csr_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  reg_csr_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  reg_csr_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  reg_csr_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  reg_csr_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  reg_csr_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  reg_csr_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  reg_csr_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  reg_csr_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  reg_csr_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  reg_csr_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  reg_csr_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  reg_csr_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  reg_csr_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  reg_csr_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  reg_csr_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  reg_csr_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  reg_csr_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  reg_csr_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  reg_csr_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  reg_csr_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  reg_csr_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  reg_csr_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  reg_csr_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  reg_csr_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  reg_csr_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  reg_csr_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  reg_csr_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  reg_csr_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  reg_csr_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  reg_csr_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  reg_csr_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  reg_csr_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  reg_csr_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  reg_csr_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  reg_csr_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  reg_csr_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  reg_csr_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  reg_csr_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  reg_csr_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  reg_csr_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  reg_csr_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  reg_csr_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  reg_csr_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  reg_csr_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  reg_csr_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  reg_csr_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  reg_csr_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  reg_csr_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  reg_csr_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  reg_csr_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  reg_csr_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  reg_csr_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  reg_csr_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  reg_csr_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  reg_csr_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  reg_csr_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  reg_csr_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  reg_csr_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  reg_csr_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  reg_csr_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  reg_csr_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  reg_csr_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  reg_csr_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  reg_csr_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  reg_csr_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  reg_csr_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  reg_csr_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  reg_csr_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  reg_csr_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  reg_csr_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  reg_csr_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  reg_csr_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  reg_csr_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  reg_csr_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  reg_csr_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  reg_csr_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  reg_csr_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  reg_csr_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  reg_csr_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  reg_csr_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  reg_csr_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  reg_csr_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  reg_csr_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  reg_csr_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  reg_csr_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  reg_csr_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  reg_csr_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  reg_csr_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  reg_csr_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  reg_csr_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  reg_csr_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  reg_csr_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  reg_csr_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  reg_csr_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  reg_csr_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  reg_csr_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  reg_csr_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  reg_csr_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  reg_csr_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  reg_csr_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  reg_csr_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  reg_csr_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  reg_csr_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  reg_csr_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  reg_csr_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  reg_csr_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  reg_csr_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  reg_csr_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  reg_csr_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  reg_csr_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  reg_csr_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  reg_csr_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  reg_csr_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  reg_csr_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  reg_csr_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  reg_csr_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  reg_csr_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  reg_csr_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  reg_csr_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  reg_csr_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  reg_csr_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  reg_csr_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  reg_csr_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  reg_csr_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  reg_csr_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  reg_csr_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  reg_csr_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  reg_csr_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  reg_csr_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  reg_csr_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  reg_csr_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  reg_csr_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  reg_csr_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  reg_csr_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  reg_csr_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  reg_csr_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  reg_csr_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  reg_csr_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  reg_csr_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  reg_csr_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  reg_csr_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  reg_csr_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  reg_csr_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  reg_csr_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  reg_csr_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  reg_csr_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  reg_csr_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  reg_csr_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  reg_csr_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  reg_csr_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  reg_csr_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  reg_csr_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  reg_csr_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  reg_csr_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  reg_csr_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  reg_csr_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  reg_csr_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  reg_csr_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  reg_csr_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  reg_csr_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  reg_csr_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  reg_csr_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  reg_csr_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  reg_csr_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  reg_csr_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  reg_csr_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  reg_csr_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  reg_csr_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  reg_csr_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  reg_csr_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  reg_csr_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  reg_csr_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  reg_csr_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  reg_csr_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  reg_csr_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  reg_csr_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  reg_csr_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  reg_csr_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  reg_csr_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  reg_csr_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  reg_csr_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  reg_csr_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  reg_csr_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  reg_csr_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  reg_csr_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  reg_csr_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  reg_csr_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  reg_csr_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  reg_csr_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  reg_csr_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  reg_csr_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  reg_csr_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  reg_csr_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  reg_csr_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  reg_csr_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  reg_csr_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  reg_csr_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  reg_csr_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  reg_csr_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  reg_csr_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  reg_csr_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  reg_csr_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  reg_csr_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  reg_csr_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  reg_csr_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  reg_csr_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  reg_csr_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  reg_csr_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  reg_csr_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  reg_csr_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  reg_csr_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  reg_csr_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  reg_csr_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  reg_csr_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  reg_csr_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  reg_csr_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  reg_csr_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  reg_csr_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  reg_csr_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  reg_csr_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  reg_csr_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  reg_csr_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  reg_csr_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  reg_csr_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  reg_csr_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  reg_csr_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  reg_csr_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  reg_csr_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  reg_csr_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  reg_csr_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  reg_csr_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  reg_csr_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  reg_csr_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  reg_csr_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  reg_csr_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  reg_csr_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  reg_csr_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  reg_csr_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  reg_csr_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  reg_csr_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  reg_csr_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  reg_csr_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  reg_csr_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  reg_csr_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  reg_csr_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  reg_csr_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  reg_csr_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  reg_csr_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  reg_csr_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  reg_csr_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  reg_csr_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  reg_csr_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  reg_csr_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  reg_csr_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  reg_csr_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  reg_csr_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  reg_csr_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  reg_csr_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  reg_csr_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  reg_csr_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  reg_csr_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  reg_csr_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  reg_csr_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  reg_csr_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  reg_csr_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  reg_csr_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  reg_csr_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  reg_csr_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  reg_csr_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  reg_csr_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  reg_csr_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  reg_csr_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  reg_csr_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  reg_csr_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  reg_csr_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  reg_csr_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  reg_csr_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  reg_csr_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  reg_csr_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  reg_csr_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  reg_csr_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  reg_csr_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  reg_csr_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  reg_csr_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  reg_csr_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  reg_csr_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  reg_csr_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  reg_csr_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  reg_csr_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  reg_csr_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  reg_csr_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  reg_csr_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  reg_csr_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  reg_csr_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  reg_csr_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  reg_csr_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  reg_csr_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  reg_csr_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  reg_csr_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  reg_csr_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  reg_csr_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  reg_csr_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  reg_csr_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  reg_csr_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  reg_csr_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  reg_csr_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  reg_csr_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  reg_csr_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  reg_csr_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  reg_csr_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  reg_csr_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  reg_csr_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  reg_csr_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  reg_csr_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  reg_csr_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  reg_csr_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  reg_csr_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  reg_csr_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  reg_csr_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  reg_csr_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  reg_csr_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  reg_csr_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  reg_csr_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  reg_csr_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  reg_csr_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  reg_csr_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  reg_csr_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  reg_csr_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  reg_csr_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  reg_csr_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  reg_csr_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  reg_csr_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  reg_csr_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  reg_csr_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  reg_csr_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  reg_csr_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  reg_csr_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  reg_csr_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  reg_csr_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  reg_csr_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  reg_csr_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  reg_csr_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  reg_csr_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  reg_csr_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  reg_csr_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  reg_csr_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  reg_csr_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  reg_csr_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  reg_csr_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  reg_csr_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  reg_csr_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  reg_csr_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  reg_csr_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  reg_csr_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  reg_csr_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  reg_csr_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  reg_csr_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  reg_csr_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  reg_csr_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  reg_csr_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  reg_csr_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  reg_csr_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  reg_csr_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  reg_csr_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  reg_csr_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  reg_csr_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  reg_csr_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  reg_csr_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  reg_csr_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  reg_csr_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  reg_csr_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  reg_csr_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  reg_csr_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  reg_csr_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  reg_csr_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  reg_csr_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  reg_csr_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  reg_csr_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  reg_csr_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  reg_csr_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  reg_csr_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  reg_csr_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  reg_csr_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  reg_csr_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  reg_csr_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  reg_csr_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  reg_csr_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  reg_csr_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  reg_csr_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  reg_csr_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  reg_csr_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  reg_csr_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  reg_csr_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  reg_csr_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  reg_csr_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  reg_csr_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  reg_csr_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  reg_csr_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  reg_csr_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  reg_csr_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  reg_csr_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  reg_csr_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  reg_csr_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  reg_csr_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  reg_csr_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  reg_csr_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  reg_csr_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  reg_csr_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  reg_csr_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  reg_csr_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  reg_csr_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  reg_csr_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  reg_csr_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  reg_csr_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  reg_csr_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  reg_csr_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  reg_csr_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  reg_csr_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  reg_csr_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  reg_csr_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  reg_csr_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  reg_csr_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  reg_csr_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  reg_csr_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  reg_csr_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  reg_csr_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  reg_csr_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  reg_csr_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  reg_csr_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  reg_csr_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  reg_csr_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  reg_csr_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  reg_csr_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  reg_csr_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  reg_csr_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  reg_csr_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  reg_csr_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  reg_csr_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  reg_csr_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  reg_csr_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  reg_csr_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  reg_csr_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  reg_csr_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  reg_csr_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  reg_csr_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  reg_csr_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  reg_csr_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  reg_csr_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  reg_csr_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  reg_csr_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  reg_csr_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  reg_csr_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  reg_csr_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  reg_csr_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  reg_csr_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  reg_csr_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  reg_csr_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  reg_csr_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  reg_csr_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  reg_csr_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  reg_csr_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  reg_csr_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  reg_csr_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  reg_csr_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  reg_csr_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  reg_csr_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  reg_csr_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  reg_csr_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  reg_csr_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  reg_csr_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  reg_csr_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  reg_csr_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  reg_csr_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  reg_csr_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  reg_csr_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  reg_csr_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  reg_csr_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  reg_csr_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  reg_csr_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  reg_csr_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  reg_csr_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  reg_csr_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  reg_csr_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  reg_csr_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  reg_csr_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  reg_csr_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  reg_csr_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  reg_csr_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  reg_csr_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  reg_csr_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  reg_csr_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  reg_csr_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  reg_csr_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  reg_csr_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  reg_csr_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  reg_csr_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  reg_csr_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  reg_csr_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  reg_csr_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  reg_csr_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  reg_csr_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  reg_csr_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  reg_csr_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  reg_csr_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  reg_csr_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  reg_csr_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  reg_csr_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  reg_csr_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  reg_csr_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  reg_csr_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  reg_csr_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  reg_csr_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  reg_csr_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  reg_csr_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  reg_csr_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  reg_csr_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  reg_csr_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  reg_csr_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  reg_csr_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  reg_csr_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  reg_csr_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  reg_csr_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  reg_csr_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  reg_csr_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  reg_csr_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  reg_csr_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  reg_csr_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  reg_csr_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  reg_csr_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  reg_csr_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  reg_csr_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  reg_csr_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  reg_csr_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  reg_csr_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  reg_csr_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  reg_csr_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  reg_csr_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  reg_csr_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  reg_csr_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  reg_csr_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  reg_csr_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  reg_csr_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  reg_csr_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  reg_csr_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  reg_csr_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  reg_csr_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  reg_csr_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  reg_csr_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  reg_csr_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  reg_csr_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  reg_csr_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  reg_csr_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  reg_csr_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  reg_csr_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  reg_csr_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  reg_csr_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  reg_csr_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  reg_csr_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  reg_csr_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  reg_csr_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  reg_csr_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  reg_csr_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  reg_csr_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  reg_csr_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  reg_csr_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  reg_csr_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  reg_csr_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  reg_csr_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  reg_csr_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  reg_csr_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  reg_csr_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  reg_csr_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  reg_csr_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  reg_csr_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  reg_csr_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  reg_csr_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  reg_csr_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  reg_csr_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  reg_csr_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  reg_csr_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  reg_csr_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  reg_csr_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  reg_csr_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  reg_csr_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  reg_csr_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  reg_csr_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  reg_csr_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  reg_csr_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  reg_csr_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  reg_csr_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  reg_csr_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  reg_csr_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  reg_csr_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  reg_csr_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  reg_csr_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  reg_csr_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  reg_csr_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  reg_csr_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  reg_csr_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  reg_csr_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  reg_csr_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  reg_csr_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  reg_csr_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  reg_csr_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  reg_csr_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  reg_csr_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  reg_csr_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  reg_csr_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  reg_csr_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  reg_csr_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  reg_csr_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  reg_csr_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  reg_csr_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  reg_csr_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  reg_csr_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  reg_csr_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  reg_csr_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  reg_csr_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  reg_csr_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  reg_csr_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  reg_csr_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  reg_csr_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  reg_csr_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  reg_csr_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  reg_csr_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  reg_csr_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  reg_csr_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  reg_csr_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  reg_csr_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  reg_csr_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  reg_csr_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  reg_csr_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  reg_csr_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  reg_csr_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  reg_csr_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  reg_csr_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  reg_csr_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  reg_csr_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  reg_csr_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  reg_csr_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  reg_csr_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  reg_csr_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  reg_csr_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  reg_csr_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  reg_csr_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  reg_csr_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  reg_csr_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  reg_csr_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  reg_csr_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  reg_csr_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  reg_csr_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  reg_csr_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  reg_csr_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  reg_csr_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  reg_csr_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  reg_csr_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  reg_csr_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  reg_csr_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  reg_csr_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  reg_csr_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  reg_csr_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  reg_csr_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  reg_csr_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  reg_csr_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  reg_csr_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  reg_csr_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  reg_csr_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  reg_csr_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  reg_csr_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  reg_csr_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  reg_csr_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  reg_csr_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  reg_csr_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  reg_csr_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  reg_csr_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  reg_csr_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  reg_csr_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  reg_csr_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  reg_csr_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  reg_csr_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  reg_csr_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  reg_csr_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  reg_csr_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  reg_csr_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  reg_csr_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  reg_csr_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  reg_csr_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  reg_csr_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  reg_csr_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  reg_csr_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  reg_csr_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  reg_csr_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  reg_csr_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  reg_csr_999 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  reg_csr_1000 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  reg_csr_1001 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  reg_csr_1002 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  reg_csr_1003 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  reg_csr_1004 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  reg_csr_1005 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  reg_csr_1006 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  reg_csr_1007 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  reg_csr_1008 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  reg_csr_1009 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  reg_csr_1010 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  reg_csr_1011 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  reg_csr_1012 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  reg_csr_1013 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  reg_csr_1014 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  reg_csr_1015 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  reg_csr_1016 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  reg_csr_1017 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  reg_csr_1018 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  reg_csr_1019 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  reg_csr_1020 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  reg_csr_1021 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  reg_csr_1022 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  reg_csr_1023 = _RAND_1023[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB(
  input         clock,
  input         reset,
  input         io_in_mem_in_rd_wen,
  input  [4:0]  io_in_mem_in_rd_addr,
  input  [31:0] io_in_mem_in_rd_data,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data
);
  wire  _T_1 = ~reset; // @[WB.scala 61:11]
  assign io_out_rd_wen = io_in_mem_in_rd_wen; // @[WB.scala 56:21]
  assign io_out_rd_addr = io_in_mem_in_rd_addr; // @[WB.scala 57:21]
  assign io_out_rd_data = io_in_mem_in_rd_data; // @[WB.scala 58:21]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------WB------------\n"); // @[WB.scala 61:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_wen: %d\n",io_in_mem_in_rd_wen); // @[WB.scala 62:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_addr: %d\n",io_in_mem_in_rd_addr); // @[WB.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_data: 0x%x\n",io_in_mem_in_rd_data); // @[WB.scala 64:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PC_BUBBLE_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_reg_pc,
  input  [31:0] io_in_inst,
  input         io_in_br_flag,
  input         io_in_jump_flag,
  input         io_stall_in_stall_flag,
  output [31:0] io_out_reg_pc,
  output [31:0] io_out_inst,
  output        io_out_br_flag,
  output        io_out_jump_flag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PC.scala 50:26]
  reg [31:0] inst; // @[PC.scala 51:26]
  wire  _inst_T = io_in_br_flag | io_in_jump_flag; // @[PC.scala 65:18]
  assign io_out_reg_pc = reg_pc; // @[PC.scala 70:25]
  assign io_out_inst = inst; // @[PC.scala 71:25]
  assign io_out_br_flag = io_in_br_flag; // @[PC.scala 72:25]
  assign io_out_jump_flag = io_in_jump_flag; // @[PC.scala 73:25]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 50:26]
      reg_pc <= 32'h0; // @[PC.scala 50:26]
    end else if (!(io_stall_in_stall_flag)) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_reg_pc;
    end
    if (reset) begin // @[PC.scala 51:26]
      inst <= 32'h0; // @[PC.scala 51:26]
    end else if (_inst_T) begin // @[Mux.scala 98:16]
      inst <= 32'h13;
    end else if (!(io_stall_in_stall_flag)) begin // @[Mux.scala 98:16]
      inst <= io_in_inst;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PC_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_reg_pc,
  output [31:0] io_out_reg_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_io_reg_reg_pc; // @[PC.scala 31:28]
  assign io_out_reg_pc = pc_io_reg_reg_pc; // @[PC.scala 34:15]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 31:28]
      pc_io_reg_reg_pc <= 32'h0; // @[PC.scala 31:28]
    end else begin
      pc_io_reg_reg_pc <= io_in_reg_pc; // @[PC.scala 33:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_io_reg_reg_pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ID_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_op1_data,
  input  [31:0] io_in_op2_data,
  input  [4:0]  io_in_rd_addr,
  input  [31:0] io_in_csr_addr_default,
  input  [4:0]  io_in_exe_fun,
  input         io_in_mem_wen,
  input         io_in_rd_wen,
  input  [2:0]  io_in_rd_sel,
  input  [2:0]  io_in_csr_cmd,
  input  [31:0] io_in_rs2_data,
  input  [31:0] io_in_imm_b_sext,
  output [31:0] io_out_op1_data,
  output [31:0] io_out_op2_data,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_csr_addr_default,
  output [4:0]  io_out_exe_fun,
  output        io_out_mem_wen,
  output        io_out_rd_wen,
  output [2:0]  io_out_rd_sel,
  output [2:0]  io_out_csr_cmd,
  output [31:0] io_out_rs2_data,
  output [31:0] io_out_imm_b_sext
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] id_io_reg_op1_data; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_op2_data; // @[ID.scala 53:28]
  reg [4:0] id_io_reg_rd_addr; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_csr_addr_default; // @[ID.scala 53:28]
  reg [4:0] id_io_reg_exe_fun; // @[ID.scala 53:28]
  reg  id_io_reg_mem_wen; // @[ID.scala 53:28]
  reg  id_io_reg_rd_wen; // @[ID.scala 53:28]
  reg [2:0] id_io_reg_rd_sel; // @[ID.scala 53:28]
  reg [2:0] id_io_reg_csr_cmd; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_rs2_data; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_imm_b_sext; // @[ID.scala 53:28]
  assign io_out_op1_data = id_io_reg_op1_data; // @[ID.scala 56:17]
  assign io_out_op2_data = id_io_reg_op2_data; // @[ID.scala 56:17]
  assign io_out_rd_addr = id_io_reg_rd_addr; // @[ID.scala 56:17]
  assign io_out_csr_addr_default = id_io_reg_csr_addr_default; // @[ID.scala 56:17]
  assign io_out_exe_fun = id_io_reg_exe_fun; // @[ID.scala 56:17]
  assign io_out_mem_wen = id_io_reg_mem_wen; // @[ID.scala 56:17]
  assign io_out_rd_wen = id_io_reg_rd_wen; // @[ID.scala 56:17]
  assign io_out_rd_sel = id_io_reg_rd_sel; // @[ID.scala 56:17]
  assign io_out_csr_cmd = id_io_reg_csr_cmd; // @[ID.scala 56:17]
  assign io_out_rs2_data = id_io_reg_rs2_data; // @[ID.scala 56:17]
  assign io_out_imm_b_sext = id_io_reg_imm_b_sext; // @[ID.scala 56:17]
  always @(posedge clock) begin
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_op1_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_op1_data <= io_in_op1_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_op2_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_op2_data <= io_in_op2_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_addr <= 5'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_addr <= io_in_rd_addr; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_csr_addr_default <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_csr_addr_default <= io_in_csr_addr_default; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_exe_fun <= 5'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_exe_fun <= io_in_exe_fun; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_mem_wen <= 1'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_mem_wen <= io_in_mem_wen; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_wen <= 1'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_wen <= io_in_rd_wen; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_sel <= 3'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_sel <= io_in_rd_sel; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_csr_cmd <= 3'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_csr_cmd <= io_in_csr_cmd; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rs2_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rs2_data <= io_in_rs2_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_imm_b_sext <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_imm_b_sext <= io_in_imm_b_sext; // @[ID.scala 55:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  id_io_reg_op1_data = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  id_io_reg_op2_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_io_reg_rd_addr = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  id_io_reg_csr_addr_default = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  id_io_reg_exe_fun = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  id_io_reg_mem_wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  id_io_reg_rd_wen = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  id_io_reg_rd_sel = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  id_io_reg_csr_cmd = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  id_io_reg_rs2_data = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  id_io_reg_imm_b_sext = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_alu_out,
  output [31:0] io_out_alu_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] alu_io_reg_alu_out; // @[ALU.scala 29:29]
  assign io_out_alu_out = alu_io_reg_alu_out; // @[ALU.scala 32:17]
  always @(posedge clock) begin
    if (reset) begin // @[ALU.scala 29:29]
      alu_io_reg_alu_out <= 32'h0; // @[ALU.scala 29:29]
    end else begin
      alu_io_reg_alu_out <= io_in_alu_out; // @[ALU.scala 31:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alu_io_reg_alu_out = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_IO_REG(
  input         clock,
  input         reset,
  input         io_in_rd_wen,
  input  [4:0]  io_in_rd_addr,
  input  [31:0] io_in_rd_data,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  wb_io_reg_rd_wen; // @[WB.scala 31:28]
  reg [4:0] wb_io_reg_rd_addr; // @[WB.scala 31:28]
  reg [31:0] wb_io_reg_rd_data; // @[WB.scala 31:28]
  assign io_out_rd_wen = wb_io_reg_rd_wen; // @[WB.scala 34:17]
  assign io_out_rd_addr = wb_io_reg_rd_addr; // @[WB.scala 34:17]
  assign io_out_rd_data = wb_io_reg_rd_data; // @[WB.scala 34:17]
  always @(posedge clock) begin
    if (reset) begin // @[WB.scala 31:28]
      wb_io_reg_rd_wen <= 1'h0; // @[WB.scala 31:28]
    end else begin
      wb_io_reg_rd_wen <= io_in_rd_wen; // @[WB.scala 33:17]
    end
    if (reset) begin // @[WB.scala 31:28]
      wb_io_reg_rd_addr <= 5'h0; // @[WB.scala 31:28]
    end else begin
      wb_io_reg_rd_addr <= io_in_rd_addr; // @[WB.scala 33:17]
    end
    if (reset) begin // @[WB.scala 31:28]
      wb_io_reg_rd_data <= 32'h0; // @[WB.scala 31:28]
    end else begin
      wb_io_reg_rd_data <= io_in_rd_data; // @[WB.scala 33:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_io_reg_rd_wen = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_io_reg_rd_addr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  wb_io_reg_rd_data = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input   clock,
  input   reset,
  output  io_exit
);
  wire  memory_clock; // @[Top.scala 15:25]
  wire [31:0] memory_io_instmem_addr; // @[Top.scala 15:25]
  wire [31:0] memory_io_instmem_inst; // @[Top.scala 15:25]
  wire [31:0] memory_io_datamem_addr; // @[Top.scala 15:25]
  wire [31:0] memory_io_datamem_rdata; // @[Top.scala 15:25]
  wire  memory_io_datamem_wen; // @[Top.scala 15:25]
  wire [31:0] memory_io_datamem_wdata; // @[Top.scala 15:25]
  wire  pc_clock; // @[Top.scala 16:25]
  wire  pc_reset; // @[Top.scala 16:25]
  wire  pc_io_in_stall_in_stall_flag; // @[Top.scala 16:25]
  wire [31:0] pc_io_in_ex_in_alu_out; // @[Top.scala 16:25]
  wire  pc_io_in_ex_in_jump_flag; // @[Top.scala 16:25]
  wire  pc_io_in_br_in_br_flag; // @[Top.scala 16:25]
  wire [31:0] pc_io_in_br_in_br_target; // @[Top.scala 16:25]
  wire [31:0] pc_io_out_reg_pc; // @[Top.scala 16:25]
  wire [31:0] pc_io_out_inst; // @[Top.scala 16:25]
  wire  pc_io_out_br_flag; // @[Top.scala 16:25]
  wire  pc_io_out_jump_flag; // @[Top.scala 16:25]
  wire [31:0] pc_io_instmem_addr; // @[Top.scala 16:25]
  wire [31:0] pc_io_instmem_inst; // @[Top.scala 16:25]
  wire  id_clock; // @[Top.scala 17:25]
  wire  id_reset; // @[Top.scala 17:25]
  wire [31:0] id_io_in_if_in_reg_pc; // @[Top.scala 17:25]
  wire [31:0] id_io_in_if_in_inst; // @[Top.scala 17:25]
  wire  id_io_in_if_in_br_flag; // @[Top.scala 17:25]
  wire  id_io_in_if_in_jump_flag; // @[Top.scala 17:25]
  wire  id_io_in_stall_in_stall_flag; // @[Top.scala 17:25]
  wire  id_io_in_mem_in_rd_wen; // @[Top.scala 17:25]
  wire [4:0] id_io_in_mem_in_rd_addr; // @[Top.scala 17:25]
  wire [31:0] id_io_in_mem_in_rd_data; // @[Top.scala 17:25]
  wire  id_io_in_wb_in_rd_wen; // @[Top.scala 17:25]
  wire [4:0] id_io_in_wb_in_rd_addr; // @[Top.scala 17:25]
  wire [31:0] id_io_in_wb_in_rd_data; // @[Top.scala 17:25]
  wire [31:0] id_io_out_op1_data; // @[Top.scala 17:25]
  wire [31:0] id_io_out_op2_data; // @[Top.scala 17:25]
  wire [4:0] id_io_out_rd_addr; // @[Top.scala 17:25]
  wire [31:0] id_io_out_csr_addr_default; // @[Top.scala 17:25]
  wire [4:0] id_io_out_exe_fun; // @[Top.scala 17:25]
  wire  id_io_out_mem_wen; // @[Top.scala 17:25]
  wire  id_io_out_rd_wen; // @[Top.scala 17:25]
  wire [2:0] id_io_out_rd_sel; // @[Top.scala 17:25]
  wire [2:0] id_io_out_csr_cmd; // @[Top.scala 17:25]
  wire [31:0] id_io_out_rs2_data; // @[Top.scala 17:25]
  wire [31:0] id_io_out_imm_b_sext; // @[Top.scala 17:25]
  wire [31:0] stall_io_in_if_in_inst; // @[Top.scala 18:25]
  wire [4:0] stall_io_in_id_reg_in_rd_addr; // @[Top.scala 18:25]
  wire  stall_io_in_id_reg_in_rd_wen; // @[Top.scala 18:25]
  wire  stall_io_out_stall_flag; // @[Top.scala 18:25]
  wire  alu_clock; // @[Top.scala 19:25]
  wire  alu_reset; // @[Top.scala 19:25]
  wire [31:0] alu_io_in_id_in_op1_data; // @[Top.scala 19:25]
  wire [31:0] alu_io_in_id_in_op2_data; // @[Top.scala 19:25]
  wire [4:0] alu_io_in_id_in_exe_fun; // @[Top.scala 19:25]
  wire [2:0] alu_io_in_id_in_rd_sel; // @[Top.scala 19:25]
  wire [31:0] alu_io_out_alu_out; // @[Top.scala 19:25]
  wire  alu_io_out_jump_flag; // @[Top.scala 19:25]
  wire  br_clock; // @[Top.scala 20:25]
  wire  br_reset; // @[Top.scala 20:25]
  wire [31:0] br_io_in_if_in_reg_pc; // @[Top.scala 20:25]
  wire [31:0] br_io_in_id_in_op1_data; // @[Top.scala 20:25]
  wire [31:0] br_io_in_id_in_op2_data; // @[Top.scala 20:25]
  wire [4:0] br_io_in_id_in_exe_fun; // @[Top.scala 20:25]
  wire [31:0] br_io_in_id_in_imm_b_sext; // @[Top.scala 20:25]
  wire  br_io_out_br_flag; // @[Top.scala 20:25]
  wire [31:0] br_io_out_br_target; // @[Top.scala 20:25]
  wire  mem_clock; // @[Top.scala 21:25]
  wire  mem_reset; // @[Top.scala 21:25]
  wire [31:0] mem_io_in_if_in_reg_pc; // @[Top.scala 21:25]
  wire [31:0] mem_io_in_id_in_op1_data; // @[Top.scala 21:25]
  wire [4:0] mem_io_in_id_in_rd_addr; // @[Top.scala 21:25]
  wire [31:0] mem_io_in_id_in_csr_addr_default; // @[Top.scala 21:25]
  wire  mem_io_in_id_in_mem_wen; // @[Top.scala 21:25]
  wire  mem_io_in_id_in_rd_wen; // @[Top.scala 21:25]
  wire [2:0] mem_io_in_id_in_rd_sel; // @[Top.scala 21:25]
  wire [2:0] mem_io_in_id_in_csr_cmd; // @[Top.scala 21:25]
  wire [31:0] mem_io_in_id_in_rs2_data; // @[Top.scala 21:25]
  wire [31:0] mem_io_in_ex_in_alu_out; // @[Top.scala 21:25]
  wire  mem_io_out_rd_wen; // @[Top.scala 21:25]
  wire [4:0] mem_io_out_rd_addr; // @[Top.scala 21:25]
  wire [31:0] mem_io_out_rd_data; // @[Top.scala 21:25]
  wire [31:0] mem_io_datamem_addr; // @[Top.scala 21:25]
  wire [31:0] mem_io_datamem_rdata; // @[Top.scala 21:25]
  wire  mem_io_datamem_wen; // @[Top.scala 21:25]
  wire [31:0] mem_io_datamem_wdata; // @[Top.scala 21:25]
  wire  wb_clock; // @[Top.scala 22:25]
  wire  wb_reset; // @[Top.scala 22:25]
  wire  wb_io_in_mem_in_rd_wen; // @[Top.scala 22:25]
  wire [4:0] wb_io_in_mem_in_rd_addr; // @[Top.scala 22:25]
  wire [31:0] wb_io_in_mem_in_rd_data; // @[Top.scala 22:25]
  wire  wb_io_out_rd_wen; // @[Top.scala 22:25]
  wire [4:0] wb_io_out_rd_addr; // @[Top.scala 22:25]
  wire [31:0] wb_io_out_rd_data; // @[Top.scala 22:25]
  wire  if_io_reg_clock; // @[Top.scala 25:33]
  wire  if_io_reg_reset; // @[Top.scala 25:33]
  wire [31:0] if_io_reg_io_in_reg_pc; // @[Top.scala 25:33]
  wire [31:0] if_io_reg_io_in_inst; // @[Top.scala 25:33]
  wire  if_io_reg_io_in_br_flag; // @[Top.scala 25:33]
  wire  if_io_reg_io_in_jump_flag; // @[Top.scala 25:33]
  wire  if_io_reg_io_stall_in_stall_flag; // @[Top.scala 25:33]
  wire [31:0] if_io_reg_io_out_reg_pc; // @[Top.scala 25:33]
  wire [31:0] if_io_reg_io_out_inst; // @[Top.scala 25:33]
  wire  if_io_reg_io_out_br_flag; // @[Top.scala 25:33]
  wire  if_io_reg_io_out_jump_flag; // @[Top.scala 25:33]
  wire  if_io_reg_n_clock; // @[Top.scala 26:33]
  wire  if_io_reg_n_reset; // @[Top.scala 26:33]
  wire [31:0] if_io_reg_n_io_in_reg_pc; // @[Top.scala 26:33]
  wire [31:0] if_io_reg_n_io_out_reg_pc; // @[Top.scala 26:33]
  wire  if_io_reg_nn_clock; // @[Top.scala 27:33]
  wire  if_io_reg_nn_reset; // @[Top.scala 27:33]
  wire [31:0] if_io_reg_nn_io_in_reg_pc; // @[Top.scala 27:33]
  wire [31:0] if_io_reg_nn_io_out_reg_pc; // @[Top.scala 27:33]
  wire  id_io_reg_clock; // @[Top.scala 28:33]
  wire  id_io_reg_reset; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_in_op1_data; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_in_op2_data; // @[Top.scala 28:33]
  wire [4:0] id_io_reg_io_in_rd_addr; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_in_csr_addr_default; // @[Top.scala 28:33]
  wire [4:0] id_io_reg_io_in_exe_fun; // @[Top.scala 28:33]
  wire  id_io_reg_io_in_mem_wen; // @[Top.scala 28:33]
  wire  id_io_reg_io_in_rd_wen; // @[Top.scala 28:33]
  wire [2:0] id_io_reg_io_in_rd_sel; // @[Top.scala 28:33]
  wire [2:0] id_io_reg_io_in_csr_cmd; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_in_rs2_data; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_in_imm_b_sext; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_out_op1_data; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_out_op2_data; // @[Top.scala 28:33]
  wire [4:0] id_io_reg_io_out_rd_addr; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_out_csr_addr_default; // @[Top.scala 28:33]
  wire [4:0] id_io_reg_io_out_exe_fun; // @[Top.scala 28:33]
  wire  id_io_reg_io_out_mem_wen; // @[Top.scala 28:33]
  wire  id_io_reg_io_out_rd_wen; // @[Top.scala 28:33]
  wire [2:0] id_io_reg_io_out_rd_sel; // @[Top.scala 28:33]
  wire [2:0] id_io_reg_io_out_csr_cmd; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_out_rs2_data; // @[Top.scala 28:33]
  wire [31:0] id_io_reg_io_out_imm_b_sext; // @[Top.scala 28:33]
  wire  id_io_reg_n_clock; // @[Top.scala 29:33]
  wire  id_io_reg_n_reset; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_in_op1_data; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_in_op2_data; // @[Top.scala 29:33]
  wire [4:0] id_io_reg_n_io_in_rd_addr; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_in_csr_addr_default; // @[Top.scala 29:33]
  wire [4:0] id_io_reg_n_io_in_exe_fun; // @[Top.scala 29:33]
  wire  id_io_reg_n_io_in_mem_wen; // @[Top.scala 29:33]
  wire  id_io_reg_n_io_in_rd_wen; // @[Top.scala 29:33]
  wire [2:0] id_io_reg_n_io_in_rd_sel; // @[Top.scala 29:33]
  wire [2:0] id_io_reg_n_io_in_csr_cmd; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_in_rs2_data; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_in_imm_b_sext; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_out_op1_data; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_out_op2_data; // @[Top.scala 29:33]
  wire [4:0] id_io_reg_n_io_out_rd_addr; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_out_csr_addr_default; // @[Top.scala 29:33]
  wire [4:0] id_io_reg_n_io_out_exe_fun; // @[Top.scala 29:33]
  wire  id_io_reg_n_io_out_mem_wen; // @[Top.scala 29:33]
  wire  id_io_reg_n_io_out_rd_wen; // @[Top.scala 29:33]
  wire [2:0] id_io_reg_n_io_out_rd_sel; // @[Top.scala 29:33]
  wire [2:0] id_io_reg_n_io_out_csr_cmd; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_out_rs2_data; // @[Top.scala 29:33]
  wire [31:0] id_io_reg_n_io_out_imm_b_sext; // @[Top.scala 29:33]
  wire  ex_io_reg_clock; // @[Top.scala 30:33]
  wire  ex_io_reg_reset; // @[Top.scala 30:33]
  wire [31:0] ex_io_reg_io_in_alu_out; // @[Top.scala 30:33]
  wire [31:0] ex_io_reg_io_out_alu_out; // @[Top.scala 30:33]
  wire  mem_io_reg_clock; // @[Top.scala 31:33]
  wire  mem_io_reg_reset; // @[Top.scala 31:33]
  wire  mem_io_reg_io_in_rd_wen; // @[Top.scala 31:33]
  wire [4:0] mem_io_reg_io_in_rd_addr; // @[Top.scala 31:33]
  wire [31:0] mem_io_reg_io_in_rd_data; // @[Top.scala 31:33]
  wire  mem_io_reg_io_out_rd_wen; // @[Top.scala 31:33]
  wire [4:0] mem_io_reg_io_out_rd_addr; // @[Top.scala 31:33]
  wire [31:0] mem_io_reg_io_out_rd_data; // @[Top.scala 31:33]
  wire [31:0] _io_exit_T = pc_io_out_inst; // @[Top.scala 79:17]
  wire  _io_exit_T_1 = 32'hc0001073 == _io_exit_T; // @[Top.scala 79:17]
  wire  _io_exit_T_2 = pc_io_out_inst == 32'h0; // @[Top.scala 80:17]
  wire  _io_exit_T_3 = pc_io_out_reg_pc == 32'h44; // @[Top.scala 81:17]
  wire  _T_1 = ~reset; // @[Top.scala 83:11]
  Memory memory ( // @[Top.scala 15:25]
    .clock(memory_clock),
    .io_instmem_addr(memory_io_instmem_addr),
    .io_instmem_inst(memory_io_instmem_inst),
    .io_datamem_addr(memory_io_datamem_addr),
    .io_datamem_rdata(memory_io_datamem_rdata),
    .io_datamem_wen(memory_io_datamem_wen),
    .io_datamem_wdata(memory_io_datamem_wdata)
  );
  PC pc ( // @[Top.scala 16:25]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_in_stall_in_stall_flag(pc_io_in_stall_in_stall_flag),
    .io_in_ex_in_alu_out(pc_io_in_ex_in_alu_out),
    .io_in_ex_in_jump_flag(pc_io_in_ex_in_jump_flag),
    .io_in_br_in_br_flag(pc_io_in_br_in_br_flag),
    .io_in_br_in_br_target(pc_io_in_br_in_br_target),
    .io_out_reg_pc(pc_io_out_reg_pc),
    .io_out_inst(pc_io_out_inst),
    .io_out_br_flag(pc_io_out_br_flag),
    .io_out_jump_flag(pc_io_out_jump_flag),
    .io_instmem_addr(pc_io_instmem_addr),
    .io_instmem_inst(pc_io_instmem_inst)
  );
  ID id ( // @[Top.scala 17:25]
    .clock(id_clock),
    .reset(id_reset),
    .io_in_if_in_reg_pc(id_io_in_if_in_reg_pc),
    .io_in_if_in_inst(id_io_in_if_in_inst),
    .io_in_if_in_br_flag(id_io_in_if_in_br_flag),
    .io_in_if_in_jump_flag(id_io_in_if_in_jump_flag),
    .io_in_stall_in_stall_flag(id_io_in_stall_in_stall_flag),
    .io_in_mem_in_rd_wen(id_io_in_mem_in_rd_wen),
    .io_in_mem_in_rd_addr(id_io_in_mem_in_rd_addr),
    .io_in_mem_in_rd_data(id_io_in_mem_in_rd_data),
    .io_in_wb_in_rd_wen(id_io_in_wb_in_rd_wen),
    .io_in_wb_in_rd_addr(id_io_in_wb_in_rd_addr),
    .io_in_wb_in_rd_data(id_io_in_wb_in_rd_data),
    .io_out_op1_data(id_io_out_op1_data),
    .io_out_op2_data(id_io_out_op2_data),
    .io_out_rd_addr(id_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_out_exe_fun),
    .io_out_mem_wen(id_io_out_mem_wen),
    .io_out_rd_wen(id_io_out_rd_wen),
    .io_out_rd_sel(id_io_out_rd_sel),
    .io_out_csr_cmd(id_io_out_csr_cmd),
    .io_out_rs2_data(id_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_out_imm_b_sext)
  );
  Stall stall ( // @[Top.scala 18:25]
    .io_in_if_in_inst(stall_io_in_if_in_inst),
    .io_in_id_reg_in_rd_addr(stall_io_in_id_reg_in_rd_addr),
    .io_in_id_reg_in_rd_wen(stall_io_in_id_reg_in_rd_wen),
    .io_out_stall_flag(stall_io_out_stall_flag)
  );
  ALU alu ( // @[Top.scala 19:25]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_id_in_op1_data(alu_io_in_id_in_op1_data),
    .io_in_id_in_op2_data(alu_io_in_id_in_op2_data),
    .io_in_id_in_exe_fun(alu_io_in_id_in_exe_fun),
    .io_in_id_in_rd_sel(alu_io_in_id_in_rd_sel),
    .io_out_alu_out(alu_io_out_alu_out),
    .io_out_jump_flag(alu_io_out_jump_flag)
  );
  BR br ( // @[Top.scala 20:25]
    .clock(br_clock),
    .reset(br_reset),
    .io_in_if_in_reg_pc(br_io_in_if_in_reg_pc),
    .io_in_id_in_op1_data(br_io_in_id_in_op1_data),
    .io_in_id_in_op2_data(br_io_in_id_in_op2_data),
    .io_in_id_in_exe_fun(br_io_in_id_in_exe_fun),
    .io_in_id_in_imm_b_sext(br_io_in_id_in_imm_b_sext),
    .io_out_br_flag(br_io_out_br_flag),
    .io_out_br_target(br_io_out_br_target)
  );
  MEM mem ( // @[Top.scala 21:25]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_if_in_reg_pc(mem_io_in_if_in_reg_pc),
    .io_in_id_in_op1_data(mem_io_in_id_in_op1_data),
    .io_in_id_in_rd_addr(mem_io_in_id_in_rd_addr),
    .io_in_id_in_csr_addr_default(mem_io_in_id_in_csr_addr_default),
    .io_in_id_in_mem_wen(mem_io_in_id_in_mem_wen),
    .io_in_id_in_rd_wen(mem_io_in_id_in_rd_wen),
    .io_in_id_in_rd_sel(mem_io_in_id_in_rd_sel),
    .io_in_id_in_csr_cmd(mem_io_in_id_in_csr_cmd),
    .io_in_id_in_rs2_data(mem_io_in_id_in_rs2_data),
    .io_in_ex_in_alu_out(mem_io_in_ex_in_alu_out),
    .io_out_rd_wen(mem_io_out_rd_wen),
    .io_out_rd_addr(mem_io_out_rd_addr),
    .io_out_rd_data(mem_io_out_rd_data),
    .io_datamem_addr(mem_io_datamem_addr),
    .io_datamem_rdata(mem_io_datamem_rdata),
    .io_datamem_wen(mem_io_datamem_wen),
    .io_datamem_wdata(mem_io_datamem_wdata)
  );
  WB wb ( // @[Top.scala 22:25]
    .clock(wb_clock),
    .reset(wb_reset),
    .io_in_mem_in_rd_wen(wb_io_in_mem_in_rd_wen),
    .io_in_mem_in_rd_addr(wb_io_in_mem_in_rd_addr),
    .io_in_mem_in_rd_data(wb_io_in_mem_in_rd_data),
    .io_out_rd_wen(wb_io_out_rd_wen),
    .io_out_rd_addr(wb_io_out_rd_addr),
    .io_out_rd_data(wb_io_out_rd_data)
  );
  PC_BUBBLE_REG if_io_reg ( // @[Top.scala 25:33]
    .clock(if_io_reg_clock),
    .reset(if_io_reg_reset),
    .io_in_reg_pc(if_io_reg_io_in_reg_pc),
    .io_in_inst(if_io_reg_io_in_inst),
    .io_in_br_flag(if_io_reg_io_in_br_flag),
    .io_in_jump_flag(if_io_reg_io_in_jump_flag),
    .io_stall_in_stall_flag(if_io_reg_io_stall_in_stall_flag),
    .io_out_reg_pc(if_io_reg_io_out_reg_pc),
    .io_out_inst(if_io_reg_io_out_inst),
    .io_out_br_flag(if_io_reg_io_out_br_flag),
    .io_out_jump_flag(if_io_reg_io_out_jump_flag)
  );
  PC_IO_REG if_io_reg_n ( // @[Top.scala 26:33]
    .clock(if_io_reg_n_clock),
    .reset(if_io_reg_n_reset),
    .io_in_reg_pc(if_io_reg_n_io_in_reg_pc),
    .io_out_reg_pc(if_io_reg_n_io_out_reg_pc)
  );
  PC_IO_REG if_io_reg_nn ( // @[Top.scala 27:33]
    .clock(if_io_reg_nn_clock),
    .reset(if_io_reg_nn_reset),
    .io_in_reg_pc(if_io_reg_nn_io_in_reg_pc),
    .io_out_reg_pc(if_io_reg_nn_io_out_reg_pc)
  );
  ID_IO_REG id_io_reg ( // @[Top.scala 28:33]
    .clock(id_io_reg_clock),
    .reset(id_io_reg_reset),
    .io_in_op1_data(id_io_reg_io_in_op1_data),
    .io_in_op2_data(id_io_reg_io_in_op2_data),
    .io_in_rd_addr(id_io_reg_io_in_rd_addr),
    .io_in_csr_addr_default(id_io_reg_io_in_csr_addr_default),
    .io_in_exe_fun(id_io_reg_io_in_exe_fun),
    .io_in_mem_wen(id_io_reg_io_in_mem_wen),
    .io_in_rd_wen(id_io_reg_io_in_rd_wen),
    .io_in_rd_sel(id_io_reg_io_in_rd_sel),
    .io_in_csr_cmd(id_io_reg_io_in_csr_cmd),
    .io_in_rs2_data(id_io_reg_io_in_rs2_data),
    .io_in_imm_b_sext(id_io_reg_io_in_imm_b_sext),
    .io_out_op1_data(id_io_reg_io_out_op1_data),
    .io_out_op2_data(id_io_reg_io_out_op2_data),
    .io_out_rd_addr(id_io_reg_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_reg_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_reg_io_out_exe_fun),
    .io_out_mem_wen(id_io_reg_io_out_mem_wen),
    .io_out_rd_wen(id_io_reg_io_out_rd_wen),
    .io_out_rd_sel(id_io_reg_io_out_rd_sel),
    .io_out_csr_cmd(id_io_reg_io_out_csr_cmd),
    .io_out_rs2_data(id_io_reg_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_reg_io_out_imm_b_sext)
  );
  ID_IO_REG id_io_reg_n ( // @[Top.scala 29:33]
    .clock(id_io_reg_n_clock),
    .reset(id_io_reg_n_reset),
    .io_in_op1_data(id_io_reg_n_io_in_op1_data),
    .io_in_op2_data(id_io_reg_n_io_in_op2_data),
    .io_in_rd_addr(id_io_reg_n_io_in_rd_addr),
    .io_in_csr_addr_default(id_io_reg_n_io_in_csr_addr_default),
    .io_in_exe_fun(id_io_reg_n_io_in_exe_fun),
    .io_in_mem_wen(id_io_reg_n_io_in_mem_wen),
    .io_in_rd_wen(id_io_reg_n_io_in_rd_wen),
    .io_in_rd_sel(id_io_reg_n_io_in_rd_sel),
    .io_in_csr_cmd(id_io_reg_n_io_in_csr_cmd),
    .io_in_rs2_data(id_io_reg_n_io_in_rs2_data),
    .io_in_imm_b_sext(id_io_reg_n_io_in_imm_b_sext),
    .io_out_op1_data(id_io_reg_n_io_out_op1_data),
    .io_out_op2_data(id_io_reg_n_io_out_op2_data),
    .io_out_rd_addr(id_io_reg_n_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_reg_n_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_reg_n_io_out_exe_fun),
    .io_out_mem_wen(id_io_reg_n_io_out_mem_wen),
    .io_out_rd_wen(id_io_reg_n_io_out_rd_wen),
    .io_out_rd_sel(id_io_reg_n_io_out_rd_sel),
    .io_out_csr_cmd(id_io_reg_n_io_out_csr_cmd),
    .io_out_rs2_data(id_io_reg_n_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_reg_n_io_out_imm_b_sext)
  );
  ALU_IO_REG ex_io_reg ( // @[Top.scala 30:33]
    .clock(ex_io_reg_clock),
    .reset(ex_io_reg_reset),
    .io_in_alu_out(ex_io_reg_io_in_alu_out),
    .io_out_alu_out(ex_io_reg_io_out_alu_out)
  );
  WB_IO_REG mem_io_reg ( // @[Top.scala 31:33]
    .clock(mem_io_reg_clock),
    .reset(mem_io_reg_reset),
    .io_in_rd_wen(mem_io_reg_io_in_rd_wen),
    .io_in_rd_addr(mem_io_reg_io_in_rd_addr),
    .io_in_rd_data(mem_io_reg_io_in_rd_data),
    .io_out_rd_wen(mem_io_reg_io_out_rd_wen),
    .io_out_rd_addr(mem_io_reg_io_out_rd_addr),
    .io_out_rd_data(mem_io_reg_io_out_rd_data)
  );
  assign io_exit = _io_exit_T_1 | (_io_exit_T_2 | _io_exit_T_3); // @[Mux.scala 98:16]
  assign memory_clock = clock;
  assign memory_io_instmem_addr = pc_io_instmem_addr; // @[Top.scala 38:25]
  assign memory_io_datamem_addr = mem_io_datamem_addr; // @[Top.scala 71:25]
  assign memory_io_datamem_wen = mem_io_datamem_wen; // @[Top.scala 71:25]
  assign memory_io_datamem_wdata = mem_io_datamem_wdata; // @[Top.scala 71:25]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_in_stall_in_stall_flag = stall_io_out_stall_flag; // @[Top.scala 35:25]
  assign pc_io_in_ex_in_alu_out = alu_io_out_alu_out; // @[Top.scala 36:25]
  assign pc_io_in_ex_in_jump_flag = alu_io_out_jump_flag; // @[Top.scala 36:25]
  assign pc_io_in_br_in_br_flag = br_io_out_br_flag; // @[Top.scala 37:25]
  assign pc_io_in_br_in_br_target = br_io_out_br_target; // @[Top.scala 37:25]
  assign pc_io_instmem_inst = memory_io_instmem_inst; // @[Top.scala 38:25]
  assign id_clock = clock;
  assign id_reset = reset;
  assign id_io_in_if_in_reg_pc = if_io_reg_io_out_reg_pc; // @[Top.scala 47:25]
  assign id_io_in_if_in_inst = if_io_reg_io_out_inst; // @[Top.scala 47:25]
  assign id_io_in_if_in_br_flag = if_io_reg_io_out_br_flag; // @[Top.scala 47:25]
  assign id_io_in_if_in_jump_flag = if_io_reg_io_out_jump_flag; // @[Top.scala 47:25]
  assign id_io_in_stall_in_stall_flag = stall_io_out_stall_flag; // @[Top.scala 49:25]
  assign id_io_in_mem_in_rd_wen = mem_io_out_rd_wen; // @[Top.scala 51:25]
  assign id_io_in_mem_in_rd_addr = mem_io_out_rd_addr; // @[Top.scala 51:25]
  assign id_io_in_mem_in_rd_data = mem_io_out_rd_data; // @[Top.scala 51:25]
  assign id_io_in_wb_in_rd_wen = wb_io_out_rd_wen; // @[Top.scala 50:25]
  assign id_io_in_wb_in_rd_addr = wb_io_out_rd_addr; // @[Top.scala 50:25]
  assign id_io_in_wb_in_rd_data = wb_io_out_rd_data; // @[Top.scala 50:25]
  assign stall_io_in_if_in_inst = if_io_reg_io_out_inst; // @[Top.scala 40:25]
  assign stall_io_in_id_reg_in_rd_addr = id_io_reg_io_out_rd_addr; // @[Top.scala 42:29]
  assign stall_io_in_id_reg_in_rd_wen = id_io_reg_io_out_rd_wen; // @[Top.scala 42:29]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_id_in_op1_data = id_io_reg_io_out_op1_data; // @[Top.scala 53:25]
  assign alu_io_in_id_in_op2_data = id_io_reg_io_out_op2_data; // @[Top.scala 53:25]
  assign alu_io_in_id_in_exe_fun = id_io_reg_io_out_exe_fun; // @[Top.scala 53:25]
  assign alu_io_in_id_in_rd_sel = id_io_reg_io_out_rd_sel; // @[Top.scala 53:25]
  assign br_clock = clock;
  assign br_reset = reset;
  assign br_io_in_if_in_reg_pc = if_io_reg_n_io_out_reg_pc; // @[Top.scala 56:25]
  assign br_io_in_id_in_op1_data = id_io_reg_io_out_op1_data; // @[Top.scala 59:25]
  assign br_io_in_id_in_op2_data = id_io_reg_io_out_op2_data; // @[Top.scala 59:25]
  assign br_io_in_id_in_exe_fun = id_io_reg_io_out_exe_fun; // @[Top.scala 59:25]
  assign br_io_in_id_in_imm_b_sext = id_io_reg_io_out_imm_b_sext; // @[Top.scala 59:25]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_if_in_reg_pc = if_io_reg_nn_io_out_reg_pc; // @[Top.scala 62:25]
  assign mem_io_in_id_in_op1_data = id_io_reg_n_io_out_op1_data; // @[Top.scala 66:25]
  assign mem_io_in_id_in_rd_addr = id_io_reg_n_io_out_rd_addr; // @[Top.scala 66:25]
  assign mem_io_in_id_in_csr_addr_default = id_io_reg_n_io_out_csr_addr_default; // @[Top.scala 66:25]
  assign mem_io_in_id_in_mem_wen = id_io_reg_n_io_out_mem_wen; // @[Top.scala 66:25]
  assign mem_io_in_id_in_rd_wen = id_io_reg_n_io_out_rd_wen; // @[Top.scala 66:25]
  assign mem_io_in_id_in_rd_sel = id_io_reg_n_io_out_rd_sel; // @[Top.scala 66:25]
  assign mem_io_in_id_in_csr_cmd = id_io_reg_n_io_out_csr_cmd; // @[Top.scala 66:25]
  assign mem_io_in_id_in_rs2_data = id_io_reg_n_io_out_rs2_data; // @[Top.scala 66:25]
  assign mem_io_in_ex_in_alu_out = ex_io_reg_io_out_alu_out; // @[Top.scala 69:25]
  assign mem_io_datamem_rdata = memory_io_datamem_rdata; // @[Top.scala 71:25]
  assign wb_clock = clock;
  assign wb_reset = reset;
  assign wb_io_in_mem_in_rd_wen = mem_io_reg_io_out_rd_wen; // @[Top.scala 73:25]
  assign wb_io_in_mem_in_rd_addr = mem_io_reg_io_out_rd_addr; // @[Top.scala 73:25]
  assign wb_io_in_mem_in_rd_data = mem_io_reg_io_out_rd_data; // @[Top.scala 73:25]
  assign if_io_reg_clock = clock;
  assign if_io_reg_reset = reset;
  assign if_io_reg_io_in_reg_pc = pc_io_out_reg_pc; // @[Top.scala 65:29]
  assign if_io_reg_io_in_inst = pc_io_out_inst; // @[Top.scala 65:29]
  assign if_io_reg_io_in_br_flag = pc_io_out_br_flag; // @[Top.scala 65:29]
  assign if_io_reg_io_in_jump_flag = pc_io_out_jump_flag; // @[Top.scala 65:29]
  assign if_io_reg_io_stall_in_stall_flag = stall_io_out_stall_flag; // @[Top.scala 45:29]
  assign if_io_reg_n_clock = clock;
  assign if_io_reg_n_reset = reset;
  assign if_io_reg_n_io_in_reg_pc = if_io_reg_io_out_reg_pc; // @[Top.scala 64:29]
  assign if_io_reg_nn_clock = clock;
  assign if_io_reg_nn_reset = reset;
  assign if_io_reg_nn_io_in_reg_pc = if_io_reg_n_io_out_reg_pc; // @[Top.scala 63:29]
  assign id_io_reg_clock = clock;
  assign id_io_reg_reset = reset;
  assign id_io_reg_io_in_op1_data = id_io_out_op1_data; // @[Top.scala 68:29]
  assign id_io_reg_io_in_op2_data = id_io_out_op2_data; // @[Top.scala 68:29]
  assign id_io_reg_io_in_rd_addr = id_io_out_rd_addr; // @[Top.scala 68:29]
  assign id_io_reg_io_in_csr_addr_default = id_io_out_csr_addr_default; // @[Top.scala 68:29]
  assign id_io_reg_io_in_exe_fun = id_io_out_exe_fun; // @[Top.scala 68:29]
  assign id_io_reg_io_in_mem_wen = id_io_out_mem_wen; // @[Top.scala 68:29]
  assign id_io_reg_io_in_rd_wen = id_io_out_rd_wen; // @[Top.scala 68:29]
  assign id_io_reg_io_in_rd_sel = id_io_out_rd_sel; // @[Top.scala 68:29]
  assign id_io_reg_io_in_csr_cmd = id_io_out_csr_cmd; // @[Top.scala 68:29]
  assign id_io_reg_io_in_rs2_data = id_io_out_rs2_data; // @[Top.scala 68:29]
  assign id_io_reg_io_in_imm_b_sext = id_io_out_imm_b_sext; // @[Top.scala 68:29]
  assign id_io_reg_n_clock = clock;
  assign id_io_reg_n_reset = reset;
  assign id_io_reg_n_io_in_op1_data = id_io_reg_io_out_op1_data; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_op2_data = id_io_reg_io_out_op2_data; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_rd_addr = id_io_reg_io_out_rd_addr; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_csr_addr_default = id_io_reg_io_out_csr_addr_default; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_exe_fun = id_io_reg_io_out_exe_fun; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_mem_wen = id_io_reg_io_out_mem_wen; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_rd_wen = id_io_reg_io_out_rd_wen; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_rd_sel = id_io_reg_io_out_rd_sel; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_csr_cmd = id_io_reg_io_out_csr_cmd; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_rs2_data = id_io_reg_io_out_rs2_data; // @[Top.scala 67:29]
  assign id_io_reg_n_io_in_imm_b_sext = id_io_reg_io_out_imm_b_sext; // @[Top.scala 67:29]
  assign ex_io_reg_clock = clock;
  assign ex_io_reg_reset = reset;
  assign ex_io_reg_io_in_alu_out = alu_io_out_alu_out; // @[Top.scala 70:29]
  assign mem_io_reg_clock = clock;
  assign mem_io_reg_reset = reset;
  assign mem_io_reg_io_in_rd_wen = mem_io_out_rd_wen; // @[Top.scala 74:29]
  assign mem_io_reg_io_in_rd_addr = mem_io_out_rd_addr; // @[Top.scala 74:29]
  assign mem_io_reg_io_in_rd_data = mem_io_out_rd_data; // @[Top.scala 74:29]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"------------------------END-----------------------\n"); // @[Top.scala 83:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"exit: %d\n",io_exit); // @[Top.scala 84:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"\n"); // @[Top.scala 85:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
