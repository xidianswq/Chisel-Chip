module Memory(
  input         clock,
  input  [31:0] io_instmem_addr,
  output [31:0] io_instmem_inst,
  input  [31:0] io_datamem_addr,
  output [31:0] io_datamem_rdata,
  input         io_datamem_wen,
  input  [31:0] io_datamem_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [7:0] mem [0:16383]; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_hi_hi_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_instmem_inst_hi_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_hi_lo_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_instmem_inst_hi_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_lo_hi_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_instmem_inst_lo_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_instmem_inst_lo_lo_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_instmem_inst_lo_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_hi_hi_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_datamem_rdata_hi_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_hi_lo_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_datamem_rdata_hi_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_lo_hi_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_datamem_rdata_lo_hi_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_io_datamem_rdata_lo_lo_data; // @[Memory.scala 45:18]
  wire [13:0] mem_io_datamem_rdata_lo_lo_addr; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_data; // @[Memory.scala 45:18]
  wire [13:0] mem_MPORT_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_1_data; // @[Memory.scala 45:18]
  wire [13:0] mem_MPORT_1_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_1_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_1_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_2_data; // @[Memory.scala 45:18]
  wire [13:0] mem_MPORT_2_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_2_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_2_en; // @[Memory.scala 45:18]
  wire [7:0] mem_MPORT_3_data; // @[Memory.scala 45:18]
  wire [13:0] mem_MPORT_3_addr; // @[Memory.scala 45:18]
  wire  mem_MPORT_3_mask; // @[Memory.scala 45:18]
  wire  mem_MPORT_3_en; // @[Memory.scala 45:18]
  wire [31:0] _io_instmem_inst_T_1 = io_instmem_addr + 32'h3; // @[Memory.scala 51:29]
  wire [31:0] _io_instmem_inst_T_4 = io_instmem_addr + 32'h2; // @[Memory.scala 52:29]
  wire [31:0] _io_instmem_inst_T_7 = io_instmem_addr + 32'h1; // @[Memory.scala 53:29]
  wire [15:0] io_instmem_inst_lo = {mem_io_instmem_inst_lo_hi_data,mem_io_instmem_inst_lo_lo_data}; // @[Cat.scala 30:58]
  wire [15:0] io_instmem_inst_hi = {mem_io_instmem_inst_hi_hi_data,mem_io_instmem_inst_hi_lo_data}; // @[Cat.scala 30:58]
  wire [31:0] _io_datamem_rdata_T_1 = io_datamem_addr + 32'h3; // @[Memory.scala 58:29]
  wire [31:0] _io_datamem_rdata_T_4 = io_datamem_addr + 32'h2; // @[Memory.scala 59:29]
  wire [31:0] _io_datamem_rdata_T_7 = io_datamem_addr + 32'h1; // @[Memory.scala 60:29]
  wire [15:0] io_datamem_rdata_lo = {mem_io_datamem_rdata_lo_hi_data,mem_io_datamem_rdata_lo_lo_data}; // @[Cat.scala 30:58]
  wire [15:0] io_datamem_rdata_hi = {mem_io_datamem_rdata_hi_hi_data,mem_io_datamem_rdata_hi_lo_data}; // @[Cat.scala 30:58]
  assign mem_io_instmem_inst_hi_hi_addr = _io_instmem_inst_T_1[13:0];
  assign mem_io_instmem_inst_hi_hi_data = mem[mem_io_instmem_inst_hi_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_hi_lo_addr = _io_instmem_inst_T_4[13:0];
  assign mem_io_instmem_inst_hi_lo_data = mem[mem_io_instmem_inst_hi_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_lo_hi_addr = _io_instmem_inst_T_7[13:0];
  assign mem_io_instmem_inst_lo_hi_data = mem[mem_io_instmem_inst_lo_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_instmem_inst_lo_lo_addr = io_instmem_addr[13:0];
  assign mem_io_instmem_inst_lo_lo_data = mem[mem_io_instmem_inst_lo_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_hi_hi_addr = _io_datamem_rdata_T_1[13:0];
  assign mem_io_datamem_rdata_hi_hi_data = mem[mem_io_datamem_rdata_hi_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_hi_lo_addr = _io_datamem_rdata_T_4[13:0];
  assign mem_io_datamem_rdata_hi_lo_data = mem[mem_io_datamem_rdata_hi_lo_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_lo_hi_addr = _io_datamem_rdata_T_7[13:0];
  assign mem_io_datamem_rdata_lo_hi_data = mem[mem_io_datamem_rdata_lo_hi_addr]; // @[Memory.scala 45:18]
  assign mem_io_datamem_rdata_lo_lo_addr = io_datamem_addr[13:0];
  assign mem_io_datamem_rdata_lo_lo_data = mem[mem_io_datamem_rdata_lo_lo_addr]; // @[Memory.scala 45:18]
  assign mem_MPORT_data = io_datamem_wdata[7:0];
  assign mem_MPORT_addr = io_datamem_addr[13:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_datamem_wen;
  assign mem_MPORT_1_data = io_datamem_wdata[15:8];
  assign mem_MPORT_1_addr = _io_datamem_rdata_T_7[13:0];
  assign mem_MPORT_1_mask = 1'h1;
  assign mem_MPORT_1_en = io_datamem_wen;
  assign mem_MPORT_2_data = io_datamem_wdata[23:16];
  assign mem_MPORT_2_addr = _io_datamem_rdata_T_4[13:0];
  assign mem_MPORT_2_mask = 1'h1;
  assign mem_MPORT_2_en = io_datamem_wen;
  assign mem_MPORT_3_data = io_datamem_wdata[31:24];
  assign mem_MPORT_3_addr = _io_datamem_rdata_T_1[13:0];
  assign mem_MPORT_3_mask = 1'h1;
  assign mem_MPORT_3_en = io_datamem_wen;
  assign io_instmem_inst = {io_instmem_inst_hi,io_instmem_inst_lo}; // @[Cat.scala 30:58]
  assign io_datamem_rdata = {io_datamem_rdata_hi,io_datamem_rdata_lo}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_1_en & mem_MPORT_1_mask) begin
      mem[mem_MPORT_1_addr] <= mem_MPORT_1_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_2_en & mem_MPORT_2_mask) begin
      mem[mem_MPORT_2_addr] <= mem_MPORT_2_data; // @[Memory.scala 45:18]
    end
    if(mem_MPORT_3_en & mem_MPORT_3_mask) begin
      mem[mem_MPORT_3_addr] <= mem_MPORT_3_data; // @[Memory.scala 45:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16384; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PC(
  input         clock,
  input         reset,
  input         io_in_bp_io_pred_flag,
  input  [31:0] io_in_bp_io_pred_target,
  input         io_in_stall_io_stall_flag,
  input         io_in_stall_io_pred_miss_flag,
  input  [31:0] io_in_ex_io_alu_io_alu_out,
  input         io_in_ex_io_alu_io_jump_flag,
  input  [31:0] io_in_ex_io_csr_io_trap_vector,
  input         io_in_ex_io_br_io_br_flag,
  input  [31:0] io_in_ex_io_br_io_br_target,
  output [31:0] io_out_reg_pc,
  output [31:0] io_out_inst,
  output [31:0] io_out_ex_io_alu_io_alu_out,
  output        io_out_ex_io_alu_io_jump_flag,
  output        io_out_ex_io_br_io_br_flag,
  output [31:0] io_out_ex_io_br_io_br_target,
  output [31:0] io_instmem_addr,
  input  [31:0] io_instmem_inst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PC.scala 104:38]
  wire [31:0] reg_pc_next_default = reg_pc + 32'h4; // @[PC.scala 105:38]
  wire  _reg_pc_next_T = io_in_stall_io_pred_miss_flag & io_in_ex_io_alu_io_jump_flag; // @[PC.scala 107:25]
  wire  _reg_pc_next_T_1 = io_in_stall_io_pred_miss_flag & io_in_ex_io_br_io_br_flag; // @[PC.scala 108:25]
  wire  _reg_pc_next_T_3 = 32'h73 == io_instmem_inst; // @[PC.scala 109:15]
  wire [31:0] _reg_pc_next_T_4 = io_in_bp_io_pred_flag ? io_in_bp_io_pred_target : reg_pc_next_default; // @[Mux.scala 98:16]
  wire [31:0] _reg_pc_next_T_5 = io_in_stall_io_stall_flag ? reg_pc : _reg_pc_next_T_4; // @[Mux.scala 98:16]
  wire  _T_1 = ~reset; // @[PC.scala 122:11]
  assign io_out_reg_pc = reg_pc; // @[PC.scala 117:25]
  assign io_out_inst = io_instmem_inst; // @[PC.scala 118:25]
  assign io_out_ex_io_alu_io_alu_out = io_in_ex_io_alu_io_alu_out; // @[PC.scala 119:25]
  assign io_out_ex_io_alu_io_jump_flag = io_in_ex_io_alu_io_jump_flag; // @[PC.scala 119:25]
  assign io_out_ex_io_br_io_br_flag = io_in_ex_io_br_io_br_flag; // @[PC.scala 119:25]
  assign io_out_ex_io_br_io_br_target = io_in_ex_io_br_io_br_target; // @[PC.scala 119:25]
  assign io_instmem_addr = reg_pc; // @[PC.scala 116:25]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 104:38]
      reg_pc <= 32'h0; // @[PC.scala 104:38]
    end else if (_reg_pc_next_T) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_ex_io_alu_io_alu_out;
    end else if (_reg_pc_next_T_1) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_ex_io_br_io_br_target;
    end else if (_reg_pc_next_T_3) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_ex_io_csr_io_trap_vector;
    end else begin
      reg_pc <= _reg_pc_next_T_5;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-----------------------START----------------------\n"); // @[PC.scala 122:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"-------------IF------------\n"); // @[PC.scala 123:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"reg_pc: 0x%x\n",reg_pc); // @[PC.scala 124:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"inst: 0x%x\n",io_instmem_inst); // @[PC.scala 125:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BP(
  input         clock,
  input         reset,
  input  [31:0] io_in_pc_io_reg_pc,
  input  [31:0] io_in_pc_io_inst,
  input  [31:0] io_in_ex_pc_io_reg_pc,
  input  [31:0] io_in_ex_io_alu_io_alu_out,
  input         io_in_ex_io_alu_io_jump_flag,
  input         io_in_ex_io_br_io_br_flag,
  input  [31:0] io_in_ex_io_br_io_br_target,
  input         io_in_ex_io_br_io_pt_flag,
  output        io_out_pred_flag,
  output [31:0] io_out_pred_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] branch_history_0; // @[BP.scala 53:42]
  reg [7:0] branch_history_1; // @[BP.scala 53:42]
  reg [7:0] branch_history_2; // @[BP.scala 53:42]
  reg [7:0] branch_history_3; // @[BP.scala 53:42]
  reg [7:0] branch_history_4; // @[BP.scala 53:42]
  reg [7:0] branch_history_5; // @[BP.scala 53:42]
  reg [7:0] branch_history_6; // @[BP.scala 53:42]
  reg [7:0] branch_history_7; // @[BP.scala 53:42]
  reg [7:0] branch_history_8; // @[BP.scala 53:42]
  reg [7:0] branch_history_9; // @[BP.scala 53:42]
  reg [7:0] branch_history_10; // @[BP.scala 53:42]
  reg [7:0] branch_history_11; // @[BP.scala 53:42]
  reg [7:0] branch_history_12; // @[BP.scala 53:42]
  reg [7:0] branch_history_13; // @[BP.scala 53:42]
  reg [7:0] branch_history_14; // @[BP.scala 53:42]
  reg [7:0] branch_history_15; // @[BP.scala 53:42]
  reg [7:0] branch_history_16; // @[BP.scala 53:42]
  reg [7:0] branch_history_17; // @[BP.scala 53:42]
  reg [7:0] branch_history_18; // @[BP.scala 53:42]
  reg [7:0] branch_history_19; // @[BP.scala 53:42]
  reg [7:0] branch_history_20; // @[BP.scala 53:42]
  reg [7:0] branch_history_21; // @[BP.scala 53:42]
  reg [7:0] branch_history_22; // @[BP.scala 53:42]
  reg [7:0] branch_history_23; // @[BP.scala 53:42]
  reg [7:0] branch_history_24; // @[BP.scala 53:42]
  reg [7:0] branch_history_25; // @[BP.scala 53:42]
  reg [7:0] branch_history_26; // @[BP.scala 53:42]
  reg [7:0] branch_history_27; // @[BP.scala 53:42]
  reg [7:0] branch_history_28; // @[BP.scala 53:42]
  reg [7:0] branch_history_29; // @[BP.scala 53:42]
  reg [7:0] branch_history_30; // @[BP.scala 53:42]
  reg [7:0] branch_history_31; // @[BP.scala 53:42]
  reg [7:0] branch_history_32; // @[BP.scala 53:42]
  reg [7:0] branch_history_33; // @[BP.scala 53:42]
  reg [7:0] branch_history_34; // @[BP.scala 53:42]
  reg [7:0] branch_history_35; // @[BP.scala 53:42]
  reg [7:0] branch_history_36; // @[BP.scala 53:42]
  reg [7:0] branch_history_37; // @[BP.scala 53:42]
  reg [7:0] branch_history_38; // @[BP.scala 53:42]
  reg [7:0] branch_history_39; // @[BP.scala 53:42]
  reg [7:0] branch_history_40; // @[BP.scala 53:42]
  reg [7:0] branch_history_41; // @[BP.scala 53:42]
  reg [7:0] branch_history_42; // @[BP.scala 53:42]
  reg [7:0] branch_history_43; // @[BP.scala 53:42]
  reg [7:0] branch_history_44; // @[BP.scala 53:42]
  reg [7:0] branch_history_45; // @[BP.scala 53:42]
  reg [7:0] branch_history_46; // @[BP.scala 53:42]
  reg [7:0] branch_history_47; // @[BP.scala 53:42]
  reg [7:0] branch_history_48; // @[BP.scala 53:42]
  reg [7:0] branch_history_49; // @[BP.scala 53:42]
  reg [7:0] branch_history_50; // @[BP.scala 53:42]
  reg [7:0] branch_history_51; // @[BP.scala 53:42]
  reg [7:0] branch_history_52; // @[BP.scala 53:42]
  reg [7:0] branch_history_53; // @[BP.scala 53:42]
  reg [7:0] branch_history_54; // @[BP.scala 53:42]
  reg [7:0] branch_history_55; // @[BP.scala 53:42]
  reg [7:0] branch_history_56; // @[BP.scala 53:42]
  reg [7:0] branch_history_57; // @[BP.scala 53:42]
  reg [7:0] branch_history_58; // @[BP.scala 53:42]
  reg [7:0] branch_history_59; // @[BP.scala 53:42]
  reg [7:0] branch_history_60; // @[BP.scala 53:42]
  reg [7:0] branch_history_61; // @[BP.scala 53:42]
  reg [7:0] branch_history_62; // @[BP.scala 53:42]
  reg [7:0] branch_history_63; // @[BP.scala 53:42]
  reg [7:0] branch_history_64; // @[BP.scala 53:42]
  reg [7:0] branch_history_65; // @[BP.scala 53:42]
  reg [7:0] branch_history_66; // @[BP.scala 53:42]
  reg [7:0] branch_history_67; // @[BP.scala 53:42]
  reg [7:0] branch_history_68; // @[BP.scala 53:42]
  reg [7:0] branch_history_69; // @[BP.scala 53:42]
  reg [7:0] branch_history_70; // @[BP.scala 53:42]
  reg [7:0] branch_history_71; // @[BP.scala 53:42]
  reg [7:0] branch_history_72; // @[BP.scala 53:42]
  reg [7:0] branch_history_73; // @[BP.scala 53:42]
  reg [7:0] branch_history_74; // @[BP.scala 53:42]
  reg [7:0] branch_history_75; // @[BP.scala 53:42]
  reg [7:0] branch_history_76; // @[BP.scala 53:42]
  reg [7:0] branch_history_77; // @[BP.scala 53:42]
  reg [7:0] branch_history_78; // @[BP.scala 53:42]
  reg [7:0] branch_history_79; // @[BP.scala 53:42]
  reg [7:0] branch_history_80; // @[BP.scala 53:42]
  reg [7:0] branch_history_81; // @[BP.scala 53:42]
  reg [7:0] branch_history_82; // @[BP.scala 53:42]
  reg [7:0] branch_history_83; // @[BP.scala 53:42]
  reg [7:0] branch_history_84; // @[BP.scala 53:42]
  reg [7:0] branch_history_85; // @[BP.scala 53:42]
  reg [7:0] branch_history_86; // @[BP.scala 53:42]
  reg [7:0] branch_history_87; // @[BP.scala 53:42]
  reg [7:0] branch_history_88; // @[BP.scala 53:42]
  reg [7:0] branch_history_89; // @[BP.scala 53:42]
  reg [7:0] branch_history_90; // @[BP.scala 53:42]
  reg [7:0] branch_history_91; // @[BP.scala 53:42]
  reg [7:0] branch_history_92; // @[BP.scala 53:42]
  reg [7:0] branch_history_93; // @[BP.scala 53:42]
  reg [7:0] branch_history_94; // @[BP.scala 53:42]
  reg [7:0] branch_history_95; // @[BP.scala 53:42]
  reg [7:0] branch_history_96; // @[BP.scala 53:42]
  reg [7:0] branch_history_97; // @[BP.scala 53:42]
  reg [7:0] branch_history_98; // @[BP.scala 53:42]
  reg [7:0] branch_history_99; // @[BP.scala 53:42]
  reg [7:0] branch_history_100; // @[BP.scala 53:42]
  reg [7:0] branch_history_101; // @[BP.scala 53:42]
  reg [7:0] branch_history_102; // @[BP.scala 53:42]
  reg [7:0] branch_history_103; // @[BP.scala 53:42]
  reg [7:0] branch_history_104; // @[BP.scala 53:42]
  reg [7:0] branch_history_105; // @[BP.scala 53:42]
  reg [7:0] branch_history_106; // @[BP.scala 53:42]
  reg [7:0] branch_history_107; // @[BP.scala 53:42]
  reg [7:0] branch_history_108; // @[BP.scala 53:42]
  reg [7:0] branch_history_109; // @[BP.scala 53:42]
  reg [7:0] branch_history_110; // @[BP.scala 53:42]
  reg [7:0] branch_history_111; // @[BP.scala 53:42]
  reg [7:0] branch_history_112; // @[BP.scala 53:42]
  reg [7:0] branch_history_113; // @[BP.scala 53:42]
  reg [7:0] branch_history_114; // @[BP.scala 53:42]
  reg [7:0] branch_history_115; // @[BP.scala 53:42]
  reg [7:0] branch_history_116; // @[BP.scala 53:42]
  reg [7:0] branch_history_117; // @[BP.scala 53:42]
  reg [7:0] branch_history_118; // @[BP.scala 53:42]
  reg [7:0] branch_history_119; // @[BP.scala 53:42]
  reg [7:0] branch_history_120; // @[BP.scala 53:42]
  reg [7:0] branch_history_121; // @[BP.scala 53:42]
  reg [7:0] branch_history_122; // @[BP.scala 53:42]
  reg [7:0] branch_history_123; // @[BP.scala 53:42]
  reg [7:0] branch_history_124; // @[BP.scala 53:42]
  reg [7:0] branch_history_125; // @[BP.scala 53:42]
  reg [7:0] branch_history_126; // @[BP.scala 53:42]
  reg [7:0] branch_history_127; // @[BP.scala 53:42]
  reg [7:0] branch_history_128; // @[BP.scala 53:42]
  reg [7:0] branch_history_129; // @[BP.scala 53:42]
  reg [7:0] branch_history_130; // @[BP.scala 53:42]
  reg [7:0] branch_history_131; // @[BP.scala 53:42]
  reg [7:0] branch_history_132; // @[BP.scala 53:42]
  reg [7:0] branch_history_133; // @[BP.scala 53:42]
  reg [7:0] branch_history_134; // @[BP.scala 53:42]
  reg [7:0] branch_history_135; // @[BP.scala 53:42]
  reg [7:0] branch_history_136; // @[BP.scala 53:42]
  reg [7:0] branch_history_137; // @[BP.scala 53:42]
  reg [7:0] branch_history_138; // @[BP.scala 53:42]
  reg [7:0] branch_history_139; // @[BP.scala 53:42]
  reg [7:0] branch_history_140; // @[BP.scala 53:42]
  reg [7:0] branch_history_141; // @[BP.scala 53:42]
  reg [7:0] branch_history_142; // @[BP.scala 53:42]
  reg [7:0] branch_history_143; // @[BP.scala 53:42]
  reg [7:0] branch_history_144; // @[BP.scala 53:42]
  reg [7:0] branch_history_145; // @[BP.scala 53:42]
  reg [7:0] branch_history_146; // @[BP.scala 53:42]
  reg [7:0] branch_history_147; // @[BP.scala 53:42]
  reg [7:0] branch_history_148; // @[BP.scala 53:42]
  reg [7:0] branch_history_149; // @[BP.scala 53:42]
  reg [7:0] branch_history_150; // @[BP.scala 53:42]
  reg [7:0] branch_history_151; // @[BP.scala 53:42]
  reg [7:0] branch_history_152; // @[BP.scala 53:42]
  reg [7:0] branch_history_153; // @[BP.scala 53:42]
  reg [7:0] branch_history_154; // @[BP.scala 53:42]
  reg [7:0] branch_history_155; // @[BP.scala 53:42]
  reg [7:0] branch_history_156; // @[BP.scala 53:42]
  reg [7:0] branch_history_157; // @[BP.scala 53:42]
  reg [7:0] branch_history_158; // @[BP.scala 53:42]
  reg [7:0] branch_history_159; // @[BP.scala 53:42]
  reg [7:0] branch_history_160; // @[BP.scala 53:42]
  reg [7:0] branch_history_161; // @[BP.scala 53:42]
  reg [7:0] branch_history_162; // @[BP.scala 53:42]
  reg [7:0] branch_history_163; // @[BP.scala 53:42]
  reg [7:0] branch_history_164; // @[BP.scala 53:42]
  reg [7:0] branch_history_165; // @[BP.scala 53:42]
  reg [7:0] branch_history_166; // @[BP.scala 53:42]
  reg [7:0] branch_history_167; // @[BP.scala 53:42]
  reg [7:0] branch_history_168; // @[BP.scala 53:42]
  reg [7:0] branch_history_169; // @[BP.scala 53:42]
  reg [7:0] branch_history_170; // @[BP.scala 53:42]
  reg [7:0] branch_history_171; // @[BP.scala 53:42]
  reg [7:0] branch_history_172; // @[BP.scala 53:42]
  reg [7:0] branch_history_173; // @[BP.scala 53:42]
  reg [7:0] branch_history_174; // @[BP.scala 53:42]
  reg [7:0] branch_history_175; // @[BP.scala 53:42]
  reg [7:0] branch_history_176; // @[BP.scala 53:42]
  reg [7:0] branch_history_177; // @[BP.scala 53:42]
  reg [7:0] branch_history_178; // @[BP.scala 53:42]
  reg [7:0] branch_history_179; // @[BP.scala 53:42]
  reg [7:0] branch_history_180; // @[BP.scala 53:42]
  reg [7:0] branch_history_181; // @[BP.scala 53:42]
  reg [7:0] branch_history_182; // @[BP.scala 53:42]
  reg [7:0] branch_history_183; // @[BP.scala 53:42]
  reg [7:0] branch_history_184; // @[BP.scala 53:42]
  reg [7:0] branch_history_185; // @[BP.scala 53:42]
  reg [7:0] branch_history_186; // @[BP.scala 53:42]
  reg [7:0] branch_history_187; // @[BP.scala 53:42]
  reg [7:0] branch_history_188; // @[BP.scala 53:42]
  reg [7:0] branch_history_189; // @[BP.scala 53:42]
  reg [7:0] branch_history_190; // @[BP.scala 53:42]
  reg [7:0] branch_history_191; // @[BP.scala 53:42]
  reg [7:0] branch_history_192; // @[BP.scala 53:42]
  reg [7:0] branch_history_193; // @[BP.scala 53:42]
  reg [7:0] branch_history_194; // @[BP.scala 53:42]
  reg [7:0] branch_history_195; // @[BP.scala 53:42]
  reg [7:0] branch_history_196; // @[BP.scala 53:42]
  reg [7:0] branch_history_197; // @[BP.scala 53:42]
  reg [7:0] branch_history_198; // @[BP.scala 53:42]
  reg [7:0] branch_history_199; // @[BP.scala 53:42]
  reg [7:0] branch_history_200; // @[BP.scala 53:42]
  reg [7:0] branch_history_201; // @[BP.scala 53:42]
  reg [7:0] branch_history_202; // @[BP.scala 53:42]
  reg [7:0] branch_history_203; // @[BP.scala 53:42]
  reg [7:0] branch_history_204; // @[BP.scala 53:42]
  reg [7:0] branch_history_205; // @[BP.scala 53:42]
  reg [7:0] branch_history_206; // @[BP.scala 53:42]
  reg [7:0] branch_history_207; // @[BP.scala 53:42]
  reg [7:0] branch_history_208; // @[BP.scala 53:42]
  reg [7:0] branch_history_209; // @[BP.scala 53:42]
  reg [7:0] branch_history_210; // @[BP.scala 53:42]
  reg [7:0] branch_history_211; // @[BP.scala 53:42]
  reg [7:0] branch_history_212; // @[BP.scala 53:42]
  reg [7:0] branch_history_213; // @[BP.scala 53:42]
  reg [7:0] branch_history_214; // @[BP.scala 53:42]
  reg [7:0] branch_history_215; // @[BP.scala 53:42]
  reg [7:0] branch_history_216; // @[BP.scala 53:42]
  reg [7:0] branch_history_217; // @[BP.scala 53:42]
  reg [7:0] branch_history_218; // @[BP.scala 53:42]
  reg [7:0] branch_history_219; // @[BP.scala 53:42]
  reg [7:0] branch_history_220; // @[BP.scala 53:42]
  reg [7:0] branch_history_221; // @[BP.scala 53:42]
  reg [7:0] branch_history_222; // @[BP.scala 53:42]
  reg [7:0] branch_history_223; // @[BP.scala 53:42]
  reg [7:0] branch_history_224; // @[BP.scala 53:42]
  reg [7:0] branch_history_225; // @[BP.scala 53:42]
  reg [7:0] branch_history_226; // @[BP.scala 53:42]
  reg [7:0] branch_history_227; // @[BP.scala 53:42]
  reg [7:0] branch_history_228; // @[BP.scala 53:42]
  reg [7:0] branch_history_229; // @[BP.scala 53:42]
  reg [7:0] branch_history_230; // @[BP.scala 53:42]
  reg [7:0] branch_history_231; // @[BP.scala 53:42]
  reg [7:0] branch_history_232; // @[BP.scala 53:42]
  reg [7:0] branch_history_233; // @[BP.scala 53:42]
  reg [7:0] branch_history_234; // @[BP.scala 53:42]
  reg [7:0] branch_history_235; // @[BP.scala 53:42]
  reg [7:0] branch_history_236; // @[BP.scala 53:42]
  reg [7:0] branch_history_237; // @[BP.scala 53:42]
  reg [7:0] branch_history_238; // @[BP.scala 53:42]
  reg [7:0] branch_history_239; // @[BP.scala 53:42]
  reg [7:0] branch_history_240; // @[BP.scala 53:42]
  reg [7:0] branch_history_241; // @[BP.scala 53:42]
  reg [7:0] branch_history_242; // @[BP.scala 53:42]
  reg [7:0] branch_history_243; // @[BP.scala 53:42]
  reg [7:0] branch_history_244; // @[BP.scala 53:42]
  reg [7:0] branch_history_245; // @[BP.scala 53:42]
  reg [7:0] branch_history_246; // @[BP.scala 53:42]
  reg [7:0] branch_history_247; // @[BP.scala 53:42]
  reg [7:0] branch_history_248; // @[BP.scala 53:42]
  reg [7:0] branch_history_249; // @[BP.scala 53:42]
  reg [7:0] branch_history_250; // @[BP.scala 53:42]
  reg [7:0] branch_history_251; // @[BP.scala 53:42]
  reg [7:0] branch_history_252; // @[BP.scala 53:42]
  reg [7:0] branch_history_253; // @[BP.scala 53:42]
  reg [7:0] branch_history_254; // @[BP.scala 53:42]
  reg [7:0] branch_history_255; // @[BP.scala 53:42]
  reg [1:0] pattern_table_0; // @[BP.scala 54:42]
  reg [1:0] pattern_table_1; // @[BP.scala 54:42]
  reg [1:0] pattern_table_2; // @[BP.scala 54:42]
  reg [1:0] pattern_table_3; // @[BP.scala 54:42]
  reg [1:0] pattern_table_4; // @[BP.scala 54:42]
  reg [1:0] pattern_table_5; // @[BP.scala 54:42]
  reg [1:0] pattern_table_6; // @[BP.scala 54:42]
  reg [1:0] pattern_table_7; // @[BP.scala 54:42]
  reg [1:0] pattern_table_8; // @[BP.scala 54:42]
  reg [1:0] pattern_table_9; // @[BP.scala 54:42]
  reg [1:0] pattern_table_10; // @[BP.scala 54:42]
  reg [1:0] pattern_table_11; // @[BP.scala 54:42]
  reg [1:0] pattern_table_12; // @[BP.scala 54:42]
  reg [1:0] pattern_table_13; // @[BP.scala 54:42]
  reg [1:0] pattern_table_14; // @[BP.scala 54:42]
  reg [1:0] pattern_table_15; // @[BP.scala 54:42]
  reg [1:0] pattern_table_16; // @[BP.scala 54:42]
  reg [1:0] pattern_table_17; // @[BP.scala 54:42]
  reg [1:0] pattern_table_18; // @[BP.scala 54:42]
  reg [1:0] pattern_table_19; // @[BP.scala 54:42]
  reg [1:0] pattern_table_20; // @[BP.scala 54:42]
  reg [1:0] pattern_table_21; // @[BP.scala 54:42]
  reg [1:0] pattern_table_22; // @[BP.scala 54:42]
  reg [1:0] pattern_table_23; // @[BP.scala 54:42]
  reg [1:0] pattern_table_24; // @[BP.scala 54:42]
  reg [1:0] pattern_table_25; // @[BP.scala 54:42]
  reg [1:0] pattern_table_26; // @[BP.scala 54:42]
  reg [1:0] pattern_table_27; // @[BP.scala 54:42]
  reg [1:0] pattern_table_28; // @[BP.scala 54:42]
  reg [1:0] pattern_table_29; // @[BP.scala 54:42]
  reg [1:0] pattern_table_30; // @[BP.scala 54:42]
  reg [1:0] pattern_table_31; // @[BP.scala 54:42]
  reg [1:0] pattern_table_32; // @[BP.scala 54:42]
  reg [1:0] pattern_table_33; // @[BP.scala 54:42]
  reg [1:0] pattern_table_34; // @[BP.scala 54:42]
  reg [1:0] pattern_table_35; // @[BP.scala 54:42]
  reg [1:0] pattern_table_36; // @[BP.scala 54:42]
  reg [1:0] pattern_table_37; // @[BP.scala 54:42]
  reg [1:0] pattern_table_38; // @[BP.scala 54:42]
  reg [1:0] pattern_table_39; // @[BP.scala 54:42]
  reg [1:0] pattern_table_40; // @[BP.scala 54:42]
  reg [1:0] pattern_table_41; // @[BP.scala 54:42]
  reg [1:0] pattern_table_42; // @[BP.scala 54:42]
  reg [1:0] pattern_table_43; // @[BP.scala 54:42]
  reg [1:0] pattern_table_44; // @[BP.scala 54:42]
  reg [1:0] pattern_table_45; // @[BP.scala 54:42]
  reg [1:0] pattern_table_46; // @[BP.scala 54:42]
  reg [1:0] pattern_table_47; // @[BP.scala 54:42]
  reg [1:0] pattern_table_48; // @[BP.scala 54:42]
  reg [1:0] pattern_table_49; // @[BP.scala 54:42]
  reg [1:0] pattern_table_50; // @[BP.scala 54:42]
  reg [1:0] pattern_table_51; // @[BP.scala 54:42]
  reg [1:0] pattern_table_52; // @[BP.scala 54:42]
  reg [1:0] pattern_table_53; // @[BP.scala 54:42]
  reg [1:0] pattern_table_54; // @[BP.scala 54:42]
  reg [1:0] pattern_table_55; // @[BP.scala 54:42]
  reg [1:0] pattern_table_56; // @[BP.scala 54:42]
  reg [1:0] pattern_table_57; // @[BP.scala 54:42]
  reg [1:0] pattern_table_58; // @[BP.scala 54:42]
  reg [1:0] pattern_table_59; // @[BP.scala 54:42]
  reg [1:0] pattern_table_60; // @[BP.scala 54:42]
  reg [1:0] pattern_table_61; // @[BP.scala 54:42]
  reg [1:0] pattern_table_62; // @[BP.scala 54:42]
  reg [1:0] pattern_table_63; // @[BP.scala 54:42]
  reg [1:0] pattern_table_64; // @[BP.scala 54:42]
  reg [1:0] pattern_table_65; // @[BP.scala 54:42]
  reg [1:0] pattern_table_66; // @[BP.scala 54:42]
  reg [1:0] pattern_table_67; // @[BP.scala 54:42]
  reg [1:0] pattern_table_68; // @[BP.scala 54:42]
  reg [1:0] pattern_table_69; // @[BP.scala 54:42]
  reg [1:0] pattern_table_70; // @[BP.scala 54:42]
  reg [1:0] pattern_table_71; // @[BP.scala 54:42]
  reg [1:0] pattern_table_72; // @[BP.scala 54:42]
  reg [1:0] pattern_table_73; // @[BP.scala 54:42]
  reg [1:0] pattern_table_74; // @[BP.scala 54:42]
  reg [1:0] pattern_table_75; // @[BP.scala 54:42]
  reg [1:0] pattern_table_76; // @[BP.scala 54:42]
  reg [1:0] pattern_table_77; // @[BP.scala 54:42]
  reg [1:0] pattern_table_78; // @[BP.scala 54:42]
  reg [1:0] pattern_table_79; // @[BP.scala 54:42]
  reg [1:0] pattern_table_80; // @[BP.scala 54:42]
  reg [1:0] pattern_table_81; // @[BP.scala 54:42]
  reg [1:0] pattern_table_82; // @[BP.scala 54:42]
  reg [1:0] pattern_table_83; // @[BP.scala 54:42]
  reg [1:0] pattern_table_84; // @[BP.scala 54:42]
  reg [1:0] pattern_table_85; // @[BP.scala 54:42]
  reg [1:0] pattern_table_86; // @[BP.scala 54:42]
  reg [1:0] pattern_table_87; // @[BP.scala 54:42]
  reg [1:0] pattern_table_88; // @[BP.scala 54:42]
  reg [1:0] pattern_table_89; // @[BP.scala 54:42]
  reg [1:0] pattern_table_90; // @[BP.scala 54:42]
  reg [1:0] pattern_table_91; // @[BP.scala 54:42]
  reg [1:0] pattern_table_92; // @[BP.scala 54:42]
  reg [1:0] pattern_table_93; // @[BP.scala 54:42]
  reg [1:0] pattern_table_94; // @[BP.scala 54:42]
  reg [1:0] pattern_table_95; // @[BP.scala 54:42]
  reg [1:0] pattern_table_96; // @[BP.scala 54:42]
  reg [1:0] pattern_table_97; // @[BP.scala 54:42]
  reg [1:0] pattern_table_98; // @[BP.scala 54:42]
  reg [1:0] pattern_table_99; // @[BP.scala 54:42]
  reg [1:0] pattern_table_100; // @[BP.scala 54:42]
  reg [1:0] pattern_table_101; // @[BP.scala 54:42]
  reg [1:0] pattern_table_102; // @[BP.scala 54:42]
  reg [1:0] pattern_table_103; // @[BP.scala 54:42]
  reg [1:0] pattern_table_104; // @[BP.scala 54:42]
  reg [1:0] pattern_table_105; // @[BP.scala 54:42]
  reg [1:0] pattern_table_106; // @[BP.scala 54:42]
  reg [1:0] pattern_table_107; // @[BP.scala 54:42]
  reg [1:0] pattern_table_108; // @[BP.scala 54:42]
  reg [1:0] pattern_table_109; // @[BP.scala 54:42]
  reg [1:0] pattern_table_110; // @[BP.scala 54:42]
  reg [1:0] pattern_table_111; // @[BP.scala 54:42]
  reg [1:0] pattern_table_112; // @[BP.scala 54:42]
  reg [1:0] pattern_table_113; // @[BP.scala 54:42]
  reg [1:0] pattern_table_114; // @[BP.scala 54:42]
  reg [1:0] pattern_table_115; // @[BP.scala 54:42]
  reg [1:0] pattern_table_116; // @[BP.scala 54:42]
  reg [1:0] pattern_table_117; // @[BP.scala 54:42]
  reg [1:0] pattern_table_118; // @[BP.scala 54:42]
  reg [1:0] pattern_table_119; // @[BP.scala 54:42]
  reg [1:0] pattern_table_120; // @[BP.scala 54:42]
  reg [1:0] pattern_table_121; // @[BP.scala 54:42]
  reg [1:0] pattern_table_122; // @[BP.scala 54:42]
  reg [1:0] pattern_table_123; // @[BP.scala 54:42]
  reg [1:0] pattern_table_124; // @[BP.scala 54:42]
  reg [1:0] pattern_table_125; // @[BP.scala 54:42]
  reg [1:0] pattern_table_126; // @[BP.scala 54:42]
  reg [1:0] pattern_table_127; // @[BP.scala 54:42]
  reg [1:0] pattern_table_128; // @[BP.scala 54:42]
  reg [1:0] pattern_table_129; // @[BP.scala 54:42]
  reg [1:0] pattern_table_130; // @[BP.scala 54:42]
  reg [1:0] pattern_table_131; // @[BP.scala 54:42]
  reg [1:0] pattern_table_132; // @[BP.scala 54:42]
  reg [1:0] pattern_table_133; // @[BP.scala 54:42]
  reg [1:0] pattern_table_134; // @[BP.scala 54:42]
  reg [1:0] pattern_table_135; // @[BP.scala 54:42]
  reg [1:0] pattern_table_136; // @[BP.scala 54:42]
  reg [1:0] pattern_table_137; // @[BP.scala 54:42]
  reg [1:0] pattern_table_138; // @[BP.scala 54:42]
  reg [1:0] pattern_table_139; // @[BP.scala 54:42]
  reg [1:0] pattern_table_140; // @[BP.scala 54:42]
  reg [1:0] pattern_table_141; // @[BP.scala 54:42]
  reg [1:0] pattern_table_142; // @[BP.scala 54:42]
  reg [1:0] pattern_table_143; // @[BP.scala 54:42]
  reg [1:0] pattern_table_144; // @[BP.scala 54:42]
  reg [1:0] pattern_table_145; // @[BP.scala 54:42]
  reg [1:0] pattern_table_146; // @[BP.scala 54:42]
  reg [1:0] pattern_table_147; // @[BP.scala 54:42]
  reg [1:0] pattern_table_148; // @[BP.scala 54:42]
  reg [1:0] pattern_table_149; // @[BP.scala 54:42]
  reg [1:0] pattern_table_150; // @[BP.scala 54:42]
  reg [1:0] pattern_table_151; // @[BP.scala 54:42]
  reg [1:0] pattern_table_152; // @[BP.scala 54:42]
  reg [1:0] pattern_table_153; // @[BP.scala 54:42]
  reg [1:0] pattern_table_154; // @[BP.scala 54:42]
  reg [1:0] pattern_table_155; // @[BP.scala 54:42]
  reg [1:0] pattern_table_156; // @[BP.scala 54:42]
  reg [1:0] pattern_table_157; // @[BP.scala 54:42]
  reg [1:0] pattern_table_158; // @[BP.scala 54:42]
  reg [1:0] pattern_table_159; // @[BP.scala 54:42]
  reg [1:0] pattern_table_160; // @[BP.scala 54:42]
  reg [1:0] pattern_table_161; // @[BP.scala 54:42]
  reg [1:0] pattern_table_162; // @[BP.scala 54:42]
  reg [1:0] pattern_table_163; // @[BP.scala 54:42]
  reg [1:0] pattern_table_164; // @[BP.scala 54:42]
  reg [1:0] pattern_table_165; // @[BP.scala 54:42]
  reg [1:0] pattern_table_166; // @[BP.scala 54:42]
  reg [1:0] pattern_table_167; // @[BP.scala 54:42]
  reg [1:0] pattern_table_168; // @[BP.scala 54:42]
  reg [1:0] pattern_table_169; // @[BP.scala 54:42]
  reg [1:0] pattern_table_170; // @[BP.scala 54:42]
  reg [1:0] pattern_table_171; // @[BP.scala 54:42]
  reg [1:0] pattern_table_172; // @[BP.scala 54:42]
  reg [1:0] pattern_table_173; // @[BP.scala 54:42]
  reg [1:0] pattern_table_174; // @[BP.scala 54:42]
  reg [1:0] pattern_table_175; // @[BP.scala 54:42]
  reg [1:0] pattern_table_176; // @[BP.scala 54:42]
  reg [1:0] pattern_table_177; // @[BP.scala 54:42]
  reg [1:0] pattern_table_178; // @[BP.scala 54:42]
  reg [1:0] pattern_table_179; // @[BP.scala 54:42]
  reg [1:0] pattern_table_180; // @[BP.scala 54:42]
  reg [1:0] pattern_table_181; // @[BP.scala 54:42]
  reg [1:0] pattern_table_182; // @[BP.scala 54:42]
  reg [1:0] pattern_table_183; // @[BP.scala 54:42]
  reg [1:0] pattern_table_184; // @[BP.scala 54:42]
  reg [1:0] pattern_table_185; // @[BP.scala 54:42]
  reg [1:0] pattern_table_186; // @[BP.scala 54:42]
  reg [1:0] pattern_table_187; // @[BP.scala 54:42]
  reg [1:0] pattern_table_188; // @[BP.scala 54:42]
  reg [1:0] pattern_table_189; // @[BP.scala 54:42]
  reg [1:0] pattern_table_190; // @[BP.scala 54:42]
  reg [1:0] pattern_table_191; // @[BP.scala 54:42]
  reg [1:0] pattern_table_192; // @[BP.scala 54:42]
  reg [1:0] pattern_table_193; // @[BP.scala 54:42]
  reg [1:0] pattern_table_194; // @[BP.scala 54:42]
  reg [1:0] pattern_table_195; // @[BP.scala 54:42]
  reg [1:0] pattern_table_196; // @[BP.scala 54:42]
  reg [1:0] pattern_table_197; // @[BP.scala 54:42]
  reg [1:0] pattern_table_198; // @[BP.scala 54:42]
  reg [1:0] pattern_table_199; // @[BP.scala 54:42]
  reg [1:0] pattern_table_200; // @[BP.scala 54:42]
  reg [1:0] pattern_table_201; // @[BP.scala 54:42]
  reg [1:0] pattern_table_202; // @[BP.scala 54:42]
  reg [1:0] pattern_table_203; // @[BP.scala 54:42]
  reg [1:0] pattern_table_204; // @[BP.scala 54:42]
  reg [1:0] pattern_table_205; // @[BP.scala 54:42]
  reg [1:0] pattern_table_206; // @[BP.scala 54:42]
  reg [1:0] pattern_table_207; // @[BP.scala 54:42]
  reg [1:0] pattern_table_208; // @[BP.scala 54:42]
  reg [1:0] pattern_table_209; // @[BP.scala 54:42]
  reg [1:0] pattern_table_210; // @[BP.scala 54:42]
  reg [1:0] pattern_table_211; // @[BP.scala 54:42]
  reg [1:0] pattern_table_212; // @[BP.scala 54:42]
  reg [1:0] pattern_table_213; // @[BP.scala 54:42]
  reg [1:0] pattern_table_214; // @[BP.scala 54:42]
  reg [1:0] pattern_table_215; // @[BP.scala 54:42]
  reg [1:0] pattern_table_216; // @[BP.scala 54:42]
  reg [1:0] pattern_table_217; // @[BP.scala 54:42]
  reg [1:0] pattern_table_218; // @[BP.scala 54:42]
  reg [1:0] pattern_table_219; // @[BP.scala 54:42]
  reg [1:0] pattern_table_220; // @[BP.scala 54:42]
  reg [1:0] pattern_table_221; // @[BP.scala 54:42]
  reg [1:0] pattern_table_222; // @[BP.scala 54:42]
  reg [1:0] pattern_table_223; // @[BP.scala 54:42]
  reg [1:0] pattern_table_224; // @[BP.scala 54:42]
  reg [1:0] pattern_table_225; // @[BP.scala 54:42]
  reg [1:0] pattern_table_226; // @[BP.scala 54:42]
  reg [1:0] pattern_table_227; // @[BP.scala 54:42]
  reg [1:0] pattern_table_228; // @[BP.scala 54:42]
  reg [1:0] pattern_table_229; // @[BP.scala 54:42]
  reg [1:0] pattern_table_230; // @[BP.scala 54:42]
  reg [1:0] pattern_table_231; // @[BP.scala 54:42]
  reg [1:0] pattern_table_232; // @[BP.scala 54:42]
  reg [1:0] pattern_table_233; // @[BP.scala 54:42]
  reg [1:0] pattern_table_234; // @[BP.scala 54:42]
  reg [1:0] pattern_table_235; // @[BP.scala 54:42]
  reg [1:0] pattern_table_236; // @[BP.scala 54:42]
  reg [1:0] pattern_table_237; // @[BP.scala 54:42]
  reg [1:0] pattern_table_238; // @[BP.scala 54:42]
  reg [1:0] pattern_table_239; // @[BP.scala 54:42]
  reg [1:0] pattern_table_240; // @[BP.scala 54:42]
  reg [1:0] pattern_table_241; // @[BP.scala 54:42]
  reg [1:0] pattern_table_242; // @[BP.scala 54:42]
  reg [1:0] pattern_table_243; // @[BP.scala 54:42]
  reg [1:0] pattern_table_244; // @[BP.scala 54:42]
  reg [1:0] pattern_table_245; // @[BP.scala 54:42]
  reg [1:0] pattern_table_246; // @[BP.scala 54:42]
  reg [1:0] pattern_table_247; // @[BP.scala 54:42]
  reg [1:0] pattern_table_248; // @[BP.scala 54:42]
  reg [1:0] pattern_table_249; // @[BP.scala 54:42]
  reg [1:0] pattern_table_250; // @[BP.scala 54:42]
  reg [1:0] pattern_table_251; // @[BP.scala 54:42]
  reg [1:0] pattern_table_252; // @[BP.scala 54:42]
  reg [1:0] pattern_table_253; // @[BP.scala 54:42]
  reg [1:0] pattern_table_254; // @[BP.scala 54:42]
  reg [1:0] pattern_table_255; // @[BP.scala 54:42]
  reg [31:0] branch_target_buffer_0; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_1; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_2; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_3; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_4; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_5; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_6; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_7; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_8; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_9; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_10; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_11; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_12; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_13; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_14; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_15; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_16; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_17; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_18; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_19; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_20; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_21; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_22; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_23; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_24; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_25; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_26; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_27; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_28; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_29; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_30; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_31; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_32; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_33; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_34; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_35; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_36; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_37; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_38; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_39; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_40; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_41; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_42; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_43; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_44; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_45; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_46; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_47; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_48; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_49; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_50; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_51; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_52; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_53; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_54; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_55; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_56; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_57; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_58; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_59; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_60; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_61; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_62; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_63; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_64; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_65; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_66; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_67; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_68; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_69; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_70; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_71; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_72; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_73; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_74; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_75; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_76; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_77; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_78; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_79; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_80; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_81; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_82; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_83; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_84; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_85; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_86; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_87; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_88; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_89; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_90; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_91; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_92; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_93; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_94; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_95; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_96; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_97; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_98; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_99; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_100; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_101; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_102; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_103; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_104; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_105; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_106; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_107; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_108; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_109; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_110; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_111; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_112; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_113; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_114; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_115; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_116; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_117; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_118; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_119; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_120; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_121; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_122; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_123; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_124; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_125; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_126; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_127; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_128; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_129; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_130; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_131; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_132; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_133; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_134; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_135; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_136; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_137; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_138; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_139; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_140; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_141; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_142; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_143; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_144; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_145; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_146; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_147; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_148; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_149; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_150; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_151; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_152; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_153; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_154; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_155; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_156; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_157; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_158; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_159; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_160; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_161; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_162; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_163; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_164; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_165; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_166; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_167; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_168; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_169; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_170; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_171; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_172; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_173; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_174; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_175; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_176; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_177; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_178; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_179; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_180; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_181; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_182; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_183; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_184; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_185; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_186; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_187; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_188; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_189; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_190; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_191; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_192; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_193; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_194; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_195; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_196; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_197; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_198; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_199; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_200; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_201; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_202; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_203; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_204; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_205; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_206; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_207; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_208; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_209; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_210; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_211; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_212; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_213; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_214; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_215; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_216; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_217; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_218; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_219; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_220; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_221; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_222; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_223; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_224; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_225; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_226; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_227; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_228; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_229; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_230; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_231; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_232; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_233; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_234; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_235; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_236; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_237; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_238; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_239; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_240; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_241; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_242; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_243; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_244; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_245; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_246; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_247; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_248; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_249; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_250; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_251; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_252; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_253; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_254; // @[BP.scala 55:42]
  reg [31:0] branch_target_buffer_255; // @[BP.scala 55:42]
  wire [7:0] ex_bh_iodex = io_in_ex_pc_io_reg_pc[9:2]; // @[BP.scala 71:32]
  wire [7:0] _GEN_1 = 8'h1 == ex_bh_iodex ? branch_history_1 : branch_history_0; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_2 = 8'h2 == ex_bh_iodex ? branch_history_2 : _GEN_1; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_3 = 8'h3 == ex_bh_iodex ? branch_history_3 : _GEN_2; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_4 = 8'h4 == ex_bh_iodex ? branch_history_4 : _GEN_3; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_5 = 8'h5 == ex_bh_iodex ? branch_history_5 : _GEN_4; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_6 = 8'h6 == ex_bh_iodex ? branch_history_6 : _GEN_5; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_7 = 8'h7 == ex_bh_iodex ? branch_history_7 : _GEN_6; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_8 = 8'h8 == ex_bh_iodex ? branch_history_8 : _GEN_7; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_9 = 8'h9 == ex_bh_iodex ? branch_history_9 : _GEN_8; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_10 = 8'ha == ex_bh_iodex ? branch_history_10 : _GEN_9; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_11 = 8'hb == ex_bh_iodex ? branch_history_11 : _GEN_10; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_12 = 8'hc == ex_bh_iodex ? branch_history_12 : _GEN_11; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_13 = 8'hd == ex_bh_iodex ? branch_history_13 : _GEN_12; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_14 = 8'he == ex_bh_iodex ? branch_history_14 : _GEN_13; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_15 = 8'hf == ex_bh_iodex ? branch_history_15 : _GEN_14; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_16 = 8'h10 == ex_bh_iodex ? branch_history_16 : _GEN_15; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_17 = 8'h11 == ex_bh_iodex ? branch_history_17 : _GEN_16; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_18 = 8'h12 == ex_bh_iodex ? branch_history_18 : _GEN_17; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_19 = 8'h13 == ex_bh_iodex ? branch_history_19 : _GEN_18; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_20 = 8'h14 == ex_bh_iodex ? branch_history_20 : _GEN_19; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_21 = 8'h15 == ex_bh_iodex ? branch_history_21 : _GEN_20; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_22 = 8'h16 == ex_bh_iodex ? branch_history_22 : _GEN_21; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_23 = 8'h17 == ex_bh_iodex ? branch_history_23 : _GEN_22; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_24 = 8'h18 == ex_bh_iodex ? branch_history_24 : _GEN_23; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_25 = 8'h19 == ex_bh_iodex ? branch_history_25 : _GEN_24; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_26 = 8'h1a == ex_bh_iodex ? branch_history_26 : _GEN_25; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_27 = 8'h1b == ex_bh_iodex ? branch_history_27 : _GEN_26; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_28 = 8'h1c == ex_bh_iodex ? branch_history_28 : _GEN_27; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_29 = 8'h1d == ex_bh_iodex ? branch_history_29 : _GEN_28; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_30 = 8'h1e == ex_bh_iodex ? branch_history_30 : _GEN_29; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_31 = 8'h1f == ex_bh_iodex ? branch_history_31 : _GEN_30; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_32 = 8'h20 == ex_bh_iodex ? branch_history_32 : _GEN_31; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_33 = 8'h21 == ex_bh_iodex ? branch_history_33 : _GEN_32; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_34 = 8'h22 == ex_bh_iodex ? branch_history_34 : _GEN_33; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_35 = 8'h23 == ex_bh_iodex ? branch_history_35 : _GEN_34; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_36 = 8'h24 == ex_bh_iodex ? branch_history_36 : _GEN_35; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_37 = 8'h25 == ex_bh_iodex ? branch_history_37 : _GEN_36; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_38 = 8'h26 == ex_bh_iodex ? branch_history_38 : _GEN_37; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_39 = 8'h27 == ex_bh_iodex ? branch_history_39 : _GEN_38; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_40 = 8'h28 == ex_bh_iodex ? branch_history_40 : _GEN_39; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_41 = 8'h29 == ex_bh_iodex ? branch_history_41 : _GEN_40; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_42 = 8'h2a == ex_bh_iodex ? branch_history_42 : _GEN_41; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_43 = 8'h2b == ex_bh_iodex ? branch_history_43 : _GEN_42; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_44 = 8'h2c == ex_bh_iodex ? branch_history_44 : _GEN_43; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_45 = 8'h2d == ex_bh_iodex ? branch_history_45 : _GEN_44; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_46 = 8'h2e == ex_bh_iodex ? branch_history_46 : _GEN_45; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_47 = 8'h2f == ex_bh_iodex ? branch_history_47 : _GEN_46; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_48 = 8'h30 == ex_bh_iodex ? branch_history_48 : _GEN_47; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_49 = 8'h31 == ex_bh_iodex ? branch_history_49 : _GEN_48; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_50 = 8'h32 == ex_bh_iodex ? branch_history_50 : _GEN_49; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_51 = 8'h33 == ex_bh_iodex ? branch_history_51 : _GEN_50; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_52 = 8'h34 == ex_bh_iodex ? branch_history_52 : _GEN_51; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_53 = 8'h35 == ex_bh_iodex ? branch_history_53 : _GEN_52; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_54 = 8'h36 == ex_bh_iodex ? branch_history_54 : _GEN_53; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_55 = 8'h37 == ex_bh_iodex ? branch_history_55 : _GEN_54; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_56 = 8'h38 == ex_bh_iodex ? branch_history_56 : _GEN_55; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_57 = 8'h39 == ex_bh_iodex ? branch_history_57 : _GEN_56; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_58 = 8'h3a == ex_bh_iodex ? branch_history_58 : _GEN_57; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_59 = 8'h3b == ex_bh_iodex ? branch_history_59 : _GEN_58; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_60 = 8'h3c == ex_bh_iodex ? branch_history_60 : _GEN_59; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_61 = 8'h3d == ex_bh_iodex ? branch_history_61 : _GEN_60; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_62 = 8'h3e == ex_bh_iodex ? branch_history_62 : _GEN_61; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_63 = 8'h3f == ex_bh_iodex ? branch_history_63 : _GEN_62; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_64 = 8'h40 == ex_bh_iodex ? branch_history_64 : _GEN_63; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_65 = 8'h41 == ex_bh_iodex ? branch_history_65 : _GEN_64; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_66 = 8'h42 == ex_bh_iodex ? branch_history_66 : _GEN_65; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_67 = 8'h43 == ex_bh_iodex ? branch_history_67 : _GEN_66; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_68 = 8'h44 == ex_bh_iodex ? branch_history_68 : _GEN_67; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_69 = 8'h45 == ex_bh_iodex ? branch_history_69 : _GEN_68; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_70 = 8'h46 == ex_bh_iodex ? branch_history_70 : _GEN_69; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_71 = 8'h47 == ex_bh_iodex ? branch_history_71 : _GEN_70; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_72 = 8'h48 == ex_bh_iodex ? branch_history_72 : _GEN_71; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_73 = 8'h49 == ex_bh_iodex ? branch_history_73 : _GEN_72; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_74 = 8'h4a == ex_bh_iodex ? branch_history_74 : _GEN_73; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_75 = 8'h4b == ex_bh_iodex ? branch_history_75 : _GEN_74; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_76 = 8'h4c == ex_bh_iodex ? branch_history_76 : _GEN_75; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_77 = 8'h4d == ex_bh_iodex ? branch_history_77 : _GEN_76; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_78 = 8'h4e == ex_bh_iodex ? branch_history_78 : _GEN_77; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_79 = 8'h4f == ex_bh_iodex ? branch_history_79 : _GEN_78; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_80 = 8'h50 == ex_bh_iodex ? branch_history_80 : _GEN_79; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_81 = 8'h51 == ex_bh_iodex ? branch_history_81 : _GEN_80; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_82 = 8'h52 == ex_bh_iodex ? branch_history_82 : _GEN_81; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_83 = 8'h53 == ex_bh_iodex ? branch_history_83 : _GEN_82; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_84 = 8'h54 == ex_bh_iodex ? branch_history_84 : _GEN_83; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_85 = 8'h55 == ex_bh_iodex ? branch_history_85 : _GEN_84; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_86 = 8'h56 == ex_bh_iodex ? branch_history_86 : _GEN_85; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_87 = 8'h57 == ex_bh_iodex ? branch_history_87 : _GEN_86; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_88 = 8'h58 == ex_bh_iodex ? branch_history_88 : _GEN_87; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_89 = 8'h59 == ex_bh_iodex ? branch_history_89 : _GEN_88; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_90 = 8'h5a == ex_bh_iodex ? branch_history_90 : _GEN_89; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_91 = 8'h5b == ex_bh_iodex ? branch_history_91 : _GEN_90; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_92 = 8'h5c == ex_bh_iodex ? branch_history_92 : _GEN_91; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_93 = 8'h5d == ex_bh_iodex ? branch_history_93 : _GEN_92; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_94 = 8'h5e == ex_bh_iodex ? branch_history_94 : _GEN_93; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_95 = 8'h5f == ex_bh_iodex ? branch_history_95 : _GEN_94; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_96 = 8'h60 == ex_bh_iodex ? branch_history_96 : _GEN_95; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_97 = 8'h61 == ex_bh_iodex ? branch_history_97 : _GEN_96; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_98 = 8'h62 == ex_bh_iodex ? branch_history_98 : _GEN_97; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_99 = 8'h63 == ex_bh_iodex ? branch_history_99 : _GEN_98; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_100 = 8'h64 == ex_bh_iodex ? branch_history_100 : _GEN_99; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_101 = 8'h65 == ex_bh_iodex ? branch_history_101 : _GEN_100; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_102 = 8'h66 == ex_bh_iodex ? branch_history_102 : _GEN_101; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_103 = 8'h67 == ex_bh_iodex ? branch_history_103 : _GEN_102; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_104 = 8'h68 == ex_bh_iodex ? branch_history_104 : _GEN_103; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_105 = 8'h69 == ex_bh_iodex ? branch_history_105 : _GEN_104; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_106 = 8'h6a == ex_bh_iodex ? branch_history_106 : _GEN_105; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_107 = 8'h6b == ex_bh_iodex ? branch_history_107 : _GEN_106; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_108 = 8'h6c == ex_bh_iodex ? branch_history_108 : _GEN_107; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_109 = 8'h6d == ex_bh_iodex ? branch_history_109 : _GEN_108; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_110 = 8'h6e == ex_bh_iodex ? branch_history_110 : _GEN_109; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_111 = 8'h6f == ex_bh_iodex ? branch_history_111 : _GEN_110; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_112 = 8'h70 == ex_bh_iodex ? branch_history_112 : _GEN_111; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_113 = 8'h71 == ex_bh_iodex ? branch_history_113 : _GEN_112; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_114 = 8'h72 == ex_bh_iodex ? branch_history_114 : _GEN_113; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_115 = 8'h73 == ex_bh_iodex ? branch_history_115 : _GEN_114; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_116 = 8'h74 == ex_bh_iodex ? branch_history_116 : _GEN_115; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_117 = 8'h75 == ex_bh_iodex ? branch_history_117 : _GEN_116; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_118 = 8'h76 == ex_bh_iodex ? branch_history_118 : _GEN_117; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_119 = 8'h77 == ex_bh_iodex ? branch_history_119 : _GEN_118; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_120 = 8'h78 == ex_bh_iodex ? branch_history_120 : _GEN_119; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_121 = 8'h79 == ex_bh_iodex ? branch_history_121 : _GEN_120; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_122 = 8'h7a == ex_bh_iodex ? branch_history_122 : _GEN_121; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_123 = 8'h7b == ex_bh_iodex ? branch_history_123 : _GEN_122; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_124 = 8'h7c == ex_bh_iodex ? branch_history_124 : _GEN_123; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_125 = 8'h7d == ex_bh_iodex ? branch_history_125 : _GEN_124; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_126 = 8'h7e == ex_bh_iodex ? branch_history_126 : _GEN_125; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_127 = 8'h7f == ex_bh_iodex ? branch_history_127 : _GEN_126; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_128 = 8'h80 == ex_bh_iodex ? branch_history_128 : _GEN_127; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_129 = 8'h81 == ex_bh_iodex ? branch_history_129 : _GEN_128; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_130 = 8'h82 == ex_bh_iodex ? branch_history_130 : _GEN_129; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_131 = 8'h83 == ex_bh_iodex ? branch_history_131 : _GEN_130; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_132 = 8'h84 == ex_bh_iodex ? branch_history_132 : _GEN_131; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_133 = 8'h85 == ex_bh_iodex ? branch_history_133 : _GEN_132; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_134 = 8'h86 == ex_bh_iodex ? branch_history_134 : _GEN_133; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_135 = 8'h87 == ex_bh_iodex ? branch_history_135 : _GEN_134; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_136 = 8'h88 == ex_bh_iodex ? branch_history_136 : _GEN_135; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_137 = 8'h89 == ex_bh_iodex ? branch_history_137 : _GEN_136; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_138 = 8'h8a == ex_bh_iodex ? branch_history_138 : _GEN_137; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_139 = 8'h8b == ex_bh_iodex ? branch_history_139 : _GEN_138; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_140 = 8'h8c == ex_bh_iodex ? branch_history_140 : _GEN_139; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_141 = 8'h8d == ex_bh_iodex ? branch_history_141 : _GEN_140; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_142 = 8'h8e == ex_bh_iodex ? branch_history_142 : _GEN_141; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_143 = 8'h8f == ex_bh_iodex ? branch_history_143 : _GEN_142; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_144 = 8'h90 == ex_bh_iodex ? branch_history_144 : _GEN_143; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_145 = 8'h91 == ex_bh_iodex ? branch_history_145 : _GEN_144; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_146 = 8'h92 == ex_bh_iodex ? branch_history_146 : _GEN_145; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_147 = 8'h93 == ex_bh_iodex ? branch_history_147 : _GEN_146; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_148 = 8'h94 == ex_bh_iodex ? branch_history_148 : _GEN_147; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_149 = 8'h95 == ex_bh_iodex ? branch_history_149 : _GEN_148; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_150 = 8'h96 == ex_bh_iodex ? branch_history_150 : _GEN_149; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_151 = 8'h97 == ex_bh_iodex ? branch_history_151 : _GEN_150; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_152 = 8'h98 == ex_bh_iodex ? branch_history_152 : _GEN_151; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_153 = 8'h99 == ex_bh_iodex ? branch_history_153 : _GEN_152; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_154 = 8'h9a == ex_bh_iodex ? branch_history_154 : _GEN_153; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_155 = 8'h9b == ex_bh_iodex ? branch_history_155 : _GEN_154; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_156 = 8'h9c == ex_bh_iodex ? branch_history_156 : _GEN_155; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_157 = 8'h9d == ex_bh_iodex ? branch_history_157 : _GEN_156; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_158 = 8'h9e == ex_bh_iodex ? branch_history_158 : _GEN_157; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_159 = 8'h9f == ex_bh_iodex ? branch_history_159 : _GEN_158; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_160 = 8'ha0 == ex_bh_iodex ? branch_history_160 : _GEN_159; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_161 = 8'ha1 == ex_bh_iodex ? branch_history_161 : _GEN_160; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_162 = 8'ha2 == ex_bh_iodex ? branch_history_162 : _GEN_161; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_163 = 8'ha3 == ex_bh_iodex ? branch_history_163 : _GEN_162; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_164 = 8'ha4 == ex_bh_iodex ? branch_history_164 : _GEN_163; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_165 = 8'ha5 == ex_bh_iodex ? branch_history_165 : _GEN_164; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_166 = 8'ha6 == ex_bh_iodex ? branch_history_166 : _GEN_165; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_167 = 8'ha7 == ex_bh_iodex ? branch_history_167 : _GEN_166; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_168 = 8'ha8 == ex_bh_iodex ? branch_history_168 : _GEN_167; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_169 = 8'ha9 == ex_bh_iodex ? branch_history_169 : _GEN_168; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_170 = 8'haa == ex_bh_iodex ? branch_history_170 : _GEN_169; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_171 = 8'hab == ex_bh_iodex ? branch_history_171 : _GEN_170; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_172 = 8'hac == ex_bh_iodex ? branch_history_172 : _GEN_171; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_173 = 8'had == ex_bh_iodex ? branch_history_173 : _GEN_172; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_174 = 8'hae == ex_bh_iodex ? branch_history_174 : _GEN_173; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_175 = 8'haf == ex_bh_iodex ? branch_history_175 : _GEN_174; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_176 = 8'hb0 == ex_bh_iodex ? branch_history_176 : _GEN_175; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_177 = 8'hb1 == ex_bh_iodex ? branch_history_177 : _GEN_176; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_178 = 8'hb2 == ex_bh_iodex ? branch_history_178 : _GEN_177; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_179 = 8'hb3 == ex_bh_iodex ? branch_history_179 : _GEN_178; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_180 = 8'hb4 == ex_bh_iodex ? branch_history_180 : _GEN_179; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_181 = 8'hb5 == ex_bh_iodex ? branch_history_181 : _GEN_180; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_182 = 8'hb6 == ex_bh_iodex ? branch_history_182 : _GEN_181; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_183 = 8'hb7 == ex_bh_iodex ? branch_history_183 : _GEN_182; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_184 = 8'hb8 == ex_bh_iodex ? branch_history_184 : _GEN_183; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_185 = 8'hb9 == ex_bh_iodex ? branch_history_185 : _GEN_184; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_186 = 8'hba == ex_bh_iodex ? branch_history_186 : _GEN_185; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_187 = 8'hbb == ex_bh_iodex ? branch_history_187 : _GEN_186; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_188 = 8'hbc == ex_bh_iodex ? branch_history_188 : _GEN_187; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_189 = 8'hbd == ex_bh_iodex ? branch_history_189 : _GEN_188; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_190 = 8'hbe == ex_bh_iodex ? branch_history_190 : _GEN_189; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_191 = 8'hbf == ex_bh_iodex ? branch_history_191 : _GEN_190; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_192 = 8'hc0 == ex_bh_iodex ? branch_history_192 : _GEN_191; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_193 = 8'hc1 == ex_bh_iodex ? branch_history_193 : _GEN_192; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_194 = 8'hc2 == ex_bh_iodex ? branch_history_194 : _GEN_193; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_195 = 8'hc3 == ex_bh_iodex ? branch_history_195 : _GEN_194; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_196 = 8'hc4 == ex_bh_iodex ? branch_history_196 : _GEN_195; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_197 = 8'hc5 == ex_bh_iodex ? branch_history_197 : _GEN_196; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_198 = 8'hc6 == ex_bh_iodex ? branch_history_198 : _GEN_197; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_199 = 8'hc7 == ex_bh_iodex ? branch_history_199 : _GEN_198; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_200 = 8'hc8 == ex_bh_iodex ? branch_history_200 : _GEN_199; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_201 = 8'hc9 == ex_bh_iodex ? branch_history_201 : _GEN_200; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_202 = 8'hca == ex_bh_iodex ? branch_history_202 : _GEN_201; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_203 = 8'hcb == ex_bh_iodex ? branch_history_203 : _GEN_202; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_204 = 8'hcc == ex_bh_iodex ? branch_history_204 : _GEN_203; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_205 = 8'hcd == ex_bh_iodex ? branch_history_205 : _GEN_204; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_206 = 8'hce == ex_bh_iodex ? branch_history_206 : _GEN_205; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_207 = 8'hcf == ex_bh_iodex ? branch_history_207 : _GEN_206; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_208 = 8'hd0 == ex_bh_iodex ? branch_history_208 : _GEN_207; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_209 = 8'hd1 == ex_bh_iodex ? branch_history_209 : _GEN_208; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_210 = 8'hd2 == ex_bh_iodex ? branch_history_210 : _GEN_209; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_211 = 8'hd3 == ex_bh_iodex ? branch_history_211 : _GEN_210; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_212 = 8'hd4 == ex_bh_iodex ? branch_history_212 : _GEN_211; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_213 = 8'hd5 == ex_bh_iodex ? branch_history_213 : _GEN_212; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_214 = 8'hd6 == ex_bh_iodex ? branch_history_214 : _GEN_213; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_215 = 8'hd7 == ex_bh_iodex ? branch_history_215 : _GEN_214; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_216 = 8'hd8 == ex_bh_iodex ? branch_history_216 : _GEN_215; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_217 = 8'hd9 == ex_bh_iodex ? branch_history_217 : _GEN_216; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_218 = 8'hda == ex_bh_iodex ? branch_history_218 : _GEN_217; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_219 = 8'hdb == ex_bh_iodex ? branch_history_219 : _GEN_218; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_220 = 8'hdc == ex_bh_iodex ? branch_history_220 : _GEN_219; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_221 = 8'hdd == ex_bh_iodex ? branch_history_221 : _GEN_220; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_222 = 8'hde == ex_bh_iodex ? branch_history_222 : _GEN_221; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_223 = 8'hdf == ex_bh_iodex ? branch_history_223 : _GEN_222; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_224 = 8'he0 == ex_bh_iodex ? branch_history_224 : _GEN_223; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_225 = 8'he1 == ex_bh_iodex ? branch_history_225 : _GEN_224; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_226 = 8'he2 == ex_bh_iodex ? branch_history_226 : _GEN_225; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_227 = 8'he3 == ex_bh_iodex ? branch_history_227 : _GEN_226; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_228 = 8'he4 == ex_bh_iodex ? branch_history_228 : _GEN_227; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_229 = 8'he5 == ex_bh_iodex ? branch_history_229 : _GEN_228; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_230 = 8'he6 == ex_bh_iodex ? branch_history_230 : _GEN_229; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_231 = 8'he7 == ex_bh_iodex ? branch_history_231 : _GEN_230; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_232 = 8'he8 == ex_bh_iodex ? branch_history_232 : _GEN_231; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_233 = 8'he9 == ex_bh_iodex ? branch_history_233 : _GEN_232; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_234 = 8'hea == ex_bh_iodex ? branch_history_234 : _GEN_233; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_235 = 8'heb == ex_bh_iodex ? branch_history_235 : _GEN_234; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_236 = 8'hec == ex_bh_iodex ? branch_history_236 : _GEN_235; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_237 = 8'hed == ex_bh_iodex ? branch_history_237 : _GEN_236; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_238 = 8'hee == ex_bh_iodex ? branch_history_238 : _GEN_237; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_239 = 8'hef == ex_bh_iodex ? branch_history_239 : _GEN_238; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_240 = 8'hf0 == ex_bh_iodex ? branch_history_240 : _GEN_239; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_241 = 8'hf1 == ex_bh_iodex ? branch_history_241 : _GEN_240; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_242 = 8'hf2 == ex_bh_iodex ? branch_history_242 : _GEN_241; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_243 = 8'hf3 == ex_bh_iodex ? branch_history_243 : _GEN_242; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_244 = 8'hf4 == ex_bh_iodex ? branch_history_244 : _GEN_243; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_245 = 8'hf5 == ex_bh_iodex ? branch_history_245 : _GEN_244; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_246 = 8'hf6 == ex_bh_iodex ? branch_history_246 : _GEN_245; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_247 = 8'hf7 == ex_bh_iodex ? branch_history_247 : _GEN_246; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_248 = 8'hf8 == ex_bh_iodex ? branch_history_248 : _GEN_247; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_249 = 8'hf9 == ex_bh_iodex ? branch_history_249 : _GEN_248; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_250 = 8'hfa == ex_bh_iodex ? branch_history_250 : _GEN_249; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_251 = 8'hfb == ex_bh_iodex ? branch_history_251 : _GEN_250; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_252 = 8'hfc == ex_bh_iodex ? branch_history_252 : _GEN_251; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_253 = 8'hfd == ex_bh_iodex ? branch_history_253 : _GEN_252; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] _GEN_254 = 8'hfe == ex_bh_iodex ? branch_history_254 : _GEN_253; // @[BP.scala 72:51 BP.scala 72:51]
  wire [7:0] ex_bh_value = 8'hff == ex_bh_iodex ? branch_history_255 : _GEN_254; // @[BP.scala 72:51 BP.scala 72:51]
  wire [8:0] _shifted_bh_T = {ex_bh_value, 1'h0}; // @[BP.scala 74:36]
  wire [7:0] shifted_bh = _shifted_bh_T[7:0]; // @[BP.scala 74:41]
  wire [7:0] _GEN_2824 = {{7'd0}, io_in_ex_io_br_io_br_flag}; // @[BP.scala 90:36]
  wire [7:0] _new_bh_value_T_2 = shifted_bh | _GEN_2824; // @[BP.scala 90:36]
  wire [7:0] new_bh_value = io_in_ex_io_br_io_pt_flag ? _new_bh_value_T_2 : shifted_bh; // @[BP.scala 88:21 BP.scala 90:22 BP.scala 87:21]
  wire [1:0] _GEN_513 = 8'h1 == ex_bh_value ? pattern_table_1 : pattern_table_0; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_514 = 8'h2 == ex_bh_value ? pattern_table_2 : _GEN_513; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_515 = 8'h3 == ex_bh_value ? pattern_table_3 : _GEN_514; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_516 = 8'h4 == ex_bh_value ? pattern_table_4 : _GEN_515; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_517 = 8'h5 == ex_bh_value ? pattern_table_5 : _GEN_516; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_518 = 8'h6 == ex_bh_value ? pattern_table_6 : _GEN_517; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_519 = 8'h7 == ex_bh_value ? pattern_table_7 : _GEN_518; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_520 = 8'h8 == ex_bh_value ? pattern_table_8 : _GEN_519; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_521 = 8'h9 == ex_bh_value ? pattern_table_9 : _GEN_520; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_522 = 8'ha == ex_bh_value ? pattern_table_10 : _GEN_521; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_523 = 8'hb == ex_bh_value ? pattern_table_11 : _GEN_522; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_524 = 8'hc == ex_bh_value ? pattern_table_12 : _GEN_523; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_525 = 8'hd == ex_bh_value ? pattern_table_13 : _GEN_524; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_526 = 8'he == ex_bh_value ? pattern_table_14 : _GEN_525; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_527 = 8'hf == ex_bh_value ? pattern_table_15 : _GEN_526; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_528 = 8'h10 == ex_bh_value ? pattern_table_16 : _GEN_527; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_529 = 8'h11 == ex_bh_value ? pattern_table_17 : _GEN_528; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_530 = 8'h12 == ex_bh_value ? pattern_table_18 : _GEN_529; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_531 = 8'h13 == ex_bh_value ? pattern_table_19 : _GEN_530; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_532 = 8'h14 == ex_bh_value ? pattern_table_20 : _GEN_531; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_533 = 8'h15 == ex_bh_value ? pattern_table_21 : _GEN_532; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_534 = 8'h16 == ex_bh_value ? pattern_table_22 : _GEN_533; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_535 = 8'h17 == ex_bh_value ? pattern_table_23 : _GEN_534; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_536 = 8'h18 == ex_bh_value ? pattern_table_24 : _GEN_535; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_537 = 8'h19 == ex_bh_value ? pattern_table_25 : _GEN_536; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_538 = 8'h1a == ex_bh_value ? pattern_table_26 : _GEN_537; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_539 = 8'h1b == ex_bh_value ? pattern_table_27 : _GEN_538; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_540 = 8'h1c == ex_bh_value ? pattern_table_28 : _GEN_539; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_541 = 8'h1d == ex_bh_value ? pattern_table_29 : _GEN_540; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_542 = 8'h1e == ex_bh_value ? pattern_table_30 : _GEN_541; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_543 = 8'h1f == ex_bh_value ? pattern_table_31 : _GEN_542; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_544 = 8'h20 == ex_bh_value ? pattern_table_32 : _GEN_543; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_545 = 8'h21 == ex_bh_value ? pattern_table_33 : _GEN_544; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_546 = 8'h22 == ex_bh_value ? pattern_table_34 : _GEN_545; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_547 = 8'h23 == ex_bh_value ? pattern_table_35 : _GEN_546; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_548 = 8'h24 == ex_bh_value ? pattern_table_36 : _GEN_547; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_549 = 8'h25 == ex_bh_value ? pattern_table_37 : _GEN_548; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_550 = 8'h26 == ex_bh_value ? pattern_table_38 : _GEN_549; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_551 = 8'h27 == ex_bh_value ? pattern_table_39 : _GEN_550; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_552 = 8'h28 == ex_bh_value ? pattern_table_40 : _GEN_551; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_553 = 8'h29 == ex_bh_value ? pattern_table_41 : _GEN_552; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_554 = 8'h2a == ex_bh_value ? pattern_table_42 : _GEN_553; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_555 = 8'h2b == ex_bh_value ? pattern_table_43 : _GEN_554; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_556 = 8'h2c == ex_bh_value ? pattern_table_44 : _GEN_555; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_557 = 8'h2d == ex_bh_value ? pattern_table_45 : _GEN_556; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_558 = 8'h2e == ex_bh_value ? pattern_table_46 : _GEN_557; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_559 = 8'h2f == ex_bh_value ? pattern_table_47 : _GEN_558; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_560 = 8'h30 == ex_bh_value ? pattern_table_48 : _GEN_559; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_561 = 8'h31 == ex_bh_value ? pattern_table_49 : _GEN_560; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_562 = 8'h32 == ex_bh_value ? pattern_table_50 : _GEN_561; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_563 = 8'h33 == ex_bh_value ? pattern_table_51 : _GEN_562; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_564 = 8'h34 == ex_bh_value ? pattern_table_52 : _GEN_563; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_565 = 8'h35 == ex_bh_value ? pattern_table_53 : _GEN_564; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_566 = 8'h36 == ex_bh_value ? pattern_table_54 : _GEN_565; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_567 = 8'h37 == ex_bh_value ? pattern_table_55 : _GEN_566; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_568 = 8'h38 == ex_bh_value ? pattern_table_56 : _GEN_567; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_569 = 8'h39 == ex_bh_value ? pattern_table_57 : _GEN_568; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_570 = 8'h3a == ex_bh_value ? pattern_table_58 : _GEN_569; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_571 = 8'h3b == ex_bh_value ? pattern_table_59 : _GEN_570; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_572 = 8'h3c == ex_bh_value ? pattern_table_60 : _GEN_571; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_573 = 8'h3d == ex_bh_value ? pattern_table_61 : _GEN_572; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_574 = 8'h3e == ex_bh_value ? pattern_table_62 : _GEN_573; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_575 = 8'h3f == ex_bh_value ? pattern_table_63 : _GEN_574; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_576 = 8'h40 == ex_bh_value ? pattern_table_64 : _GEN_575; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_577 = 8'h41 == ex_bh_value ? pattern_table_65 : _GEN_576; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_578 = 8'h42 == ex_bh_value ? pattern_table_66 : _GEN_577; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_579 = 8'h43 == ex_bh_value ? pattern_table_67 : _GEN_578; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_580 = 8'h44 == ex_bh_value ? pattern_table_68 : _GEN_579; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_581 = 8'h45 == ex_bh_value ? pattern_table_69 : _GEN_580; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_582 = 8'h46 == ex_bh_value ? pattern_table_70 : _GEN_581; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_583 = 8'h47 == ex_bh_value ? pattern_table_71 : _GEN_582; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_584 = 8'h48 == ex_bh_value ? pattern_table_72 : _GEN_583; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_585 = 8'h49 == ex_bh_value ? pattern_table_73 : _GEN_584; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_586 = 8'h4a == ex_bh_value ? pattern_table_74 : _GEN_585; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_587 = 8'h4b == ex_bh_value ? pattern_table_75 : _GEN_586; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_588 = 8'h4c == ex_bh_value ? pattern_table_76 : _GEN_587; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_589 = 8'h4d == ex_bh_value ? pattern_table_77 : _GEN_588; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_590 = 8'h4e == ex_bh_value ? pattern_table_78 : _GEN_589; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_591 = 8'h4f == ex_bh_value ? pattern_table_79 : _GEN_590; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_592 = 8'h50 == ex_bh_value ? pattern_table_80 : _GEN_591; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_593 = 8'h51 == ex_bh_value ? pattern_table_81 : _GEN_592; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_594 = 8'h52 == ex_bh_value ? pattern_table_82 : _GEN_593; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_595 = 8'h53 == ex_bh_value ? pattern_table_83 : _GEN_594; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_596 = 8'h54 == ex_bh_value ? pattern_table_84 : _GEN_595; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_597 = 8'h55 == ex_bh_value ? pattern_table_85 : _GEN_596; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_598 = 8'h56 == ex_bh_value ? pattern_table_86 : _GEN_597; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_599 = 8'h57 == ex_bh_value ? pattern_table_87 : _GEN_598; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_600 = 8'h58 == ex_bh_value ? pattern_table_88 : _GEN_599; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_601 = 8'h59 == ex_bh_value ? pattern_table_89 : _GEN_600; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_602 = 8'h5a == ex_bh_value ? pattern_table_90 : _GEN_601; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_603 = 8'h5b == ex_bh_value ? pattern_table_91 : _GEN_602; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_604 = 8'h5c == ex_bh_value ? pattern_table_92 : _GEN_603; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_605 = 8'h5d == ex_bh_value ? pattern_table_93 : _GEN_604; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_606 = 8'h5e == ex_bh_value ? pattern_table_94 : _GEN_605; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_607 = 8'h5f == ex_bh_value ? pattern_table_95 : _GEN_606; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_608 = 8'h60 == ex_bh_value ? pattern_table_96 : _GEN_607; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_609 = 8'h61 == ex_bh_value ? pattern_table_97 : _GEN_608; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_610 = 8'h62 == ex_bh_value ? pattern_table_98 : _GEN_609; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_611 = 8'h63 == ex_bh_value ? pattern_table_99 : _GEN_610; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_612 = 8'h64 == ex_bh_value ? pattern_table_100 : _GEN_611; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_613 = 8'h65 == ex_bh_value ? pattern_table_101 : _GEN_612; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_614 = 8'h66 == ex_bh_value ? pattern_table_102 : _GEN_613; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_615 = 8'h67 == ex_bh_value ? pattern_table_103 : _GEN_614; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_616 = 8'h68 == ex_bh_value ? pattern_table_104 : _GEN_615; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_617 = 8'h69 == ex_bh_value ? pattern_table_105 : _GEN_616; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_618 = 8'h6a == ex_bh_value ? pattern_table_106 : _GEN_617; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_619 = 8'h6b == ex_bh_value ? pattern_table_107 : _GEN_618; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_620 = 8'h6c == ex_bh_value ? pattern_table_108 : _GEN_619; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_621 = 8'h6d == ex_bh_value ? pattern_table_109 : _GEN_620; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_622 = 8'h6e == ex_bh_value ? pattern_table_110 : _GEN_621; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_623 = 8'h6f == ex_bh_value ? pattern_table_111 : _GEN_622; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_624 = 8'h70 == ex_bh_value ? pattern_table_112 : _GEN_623; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_625 = 8'h71 == ex_bh_value ? pattern_table_113 : _GEN_624; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_626 = 8'h72 == ex_bh_value ? pattern_table_114 : _GEN_625; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_627 = 8'h73 == ex_bh_value ? pattern_table_115 : _GEN_626; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_628 = 8'h74 == ex_bh_value ? pattern_table_116 : _GEN_627; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_629 = 8'h75 == ex_bh_value ? pattern_table_117 : _GEN_628; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_630 = 8'h76 == ex_bh_value ? pattern_table_118 : _GEN_629; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_631 = 8'h77 == ex_bh_value ? pattern_table_119 : _GEN_630; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_632 = 8'h78 == ex_bh_value ? pattern_table_120 : _GEN_631; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_633 = 8'h79 == ex_bh_value ? pattern_table_121 : _GEN_632; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_634 = 8'h7a == ex_bh_value ? pattern_table_122 : _GEN_633; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_635 = 8'h7b == ex_bh_value ? pattern_table_123 : _GEN_634; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_636 = 8'h7c == ex_bh_value ? pattern_table_124 : _GEN_635; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_637 = 8'h7d == ex_bh_value ? pattern_table_125 : _GEN_636; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_638 = 8'h7e == ex_bh_value ? pattern_table_126 : _GEN_637; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_639 = 8'h7f == ex_bh_value ? pattern_table_127 : _GEN_638; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_640 = 8'h80 == ex_bh_value ? pattern_table_128 : _GEN_639; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_641 = 8'h81 == ex_bh_value ? pattern_table_129 : _GEN_640; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_642 = 8'h82 == ex_bh_value ? pattern_table_130 : _GEN_641; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_643 = 8'h83 == ex_bh_value ? pattern_table_131 : _GEN_642; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_644 = 8'h84 == ex_bh_value ? pattern_table_132 : _GEN_643; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_645 = 8'h85 == ex_bh_value ? pattern_table_133 : _GEN_644; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_646 = 8'h86 == ex_bh_value ? pattern_table_134 : _GEN_645; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_647 = 8'h87 == ex_bh_value ? pattern_table_135 : _GEN_646; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_648 = 8'h88 == ex_bh_value ? pattern_table_136 : _GEN_647; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_649 = 8'h89 == ex_bh_value ? pattern_table_137 : _GEN_648; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_650 = 8'h8a == ex_bh_value ? pattern_table_138 : _GEN_649; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_651 = 8'h8b == ex_bh_value ? pattern_table_139 : _GEN_650; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_652 = 8'h8c == ex_bh_value ? pattern_table_140 : _GEN_651; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_653 = 8'h8d == ex_bh_value ? pattern_table_141 : _GEN_652; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_654 = 8'h8e == ex_bh_value ? pattern_table_142 : _GEN_653; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_655 = 8'h8f == ex_bh_value ? pattern_table_143 : _GEN_654; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_656 = 8'h90 == ex_bh_value ? pattern_table_144 : _GEN_655; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_657 = 8'h91 == ex_bh_value ? pattern_table_145 : _GEN_656; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_658 = 8'h92 == ex_bh_value ? pattern_table_146 : _GEN_657; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_659 = 8'h93 == ex_bh_value ? pattern_table_147 : _GEN_658; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_660 = 8'h94 == ex_bh_value ? pattern_table_148 : _GEN_659; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_661 = 8'h95 == ex_bh_value ? pattern_table_149 : _GEN_660; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_662 = 8'h96 == ex_bh_value ? pattern_table_150 : _GEN_661; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_663 = 8'h97 == ex_bh_value ? pattern_table_151 : _GEN_662; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_664 = 8'h98 == ex_bh_value ? pattern_table_152 : _GEN_663; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_665 = 8'h99 == ex_bh_value ? pattern_table_153 : _GEN_664; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_666 = 8'h9a == ex_bh_value ? pattern_table_154 : _GEN_665; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_667 = 8'h9b == ex_bh_value ? pattern_table_155 : _GEN_666; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_668 = 8'h9c == ex_bh_value ? pattern_table_156 : _GEN_667; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_669 = 8'h9d == ex_bh_value ? pattern_table_157 : _GEN_668; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_670 = 8'h9e == ex_bh_value ? pattern_table_158 : _GEN_669; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_671 = 8'h9f == ex_bh_value ? pattern_table_159 : _GEN_670; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_672 = 8'ha0 == ex_bh_value ? pattern_table_160 : _GEN_671; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_673 = 8'ha1 == ex_bh_value ? pattern_table_161 : _GEN_672; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_674 = 8'ha2 == ex_bh_value ? pattern_table_162 : _GEN_673; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_675 = 8'ha3 == ex_bh_value ? pattern_table_163 : _GEN_674; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_676 = 8'ha4 == ex_bh_value ? pattern_table_164 : _GEN_675; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_677 = 8'ha5 == ex_bh_value ? pattern_table_165 : _GEN_676; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_678 = 8'ha6 == ex_bh_value ? pattern_table_166 : _GEN_677; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_679 = 8'ha7 == ex_bh_value ? pattern_table_167 : _GEN_678; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_680 = 8'ha8 == ex_bh_value ? pattern_table_168 : _GEN_679; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_681 = 8'ha9 == ex_bh_value ? pattern_table_169 : _GEN_680; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_682 = 8'haa == ex_bh_value ? pattern_table_170 : _GEN_681; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_683 = 8'hab == ex_bh_value ? pattern_table_171 : _GEN_682; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_684 = 8'hac == ex_bh_value ? pattern_table_172 : _GEN_683; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_685 = 8'had == ex_bh_value ? pattern_table_173 : _GEN_684; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_686 = 8'hae == ex_bh_value ? pattern_table_174 : _GEN_685; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_687 = 8'haf == ex_bh_value ? pattern_table_175 : _GEN_686; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_688 = 8'hb0 == ex_bh_value ? pattern_table_176 : _GEN_687; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_689 = 8'hb1 == ex_bh_value ? pattern_table_177 : _GEN_688; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_690 = 8'hb2 == ex_bh_value ? pattern_table_178 : _GEN_689; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_691 = 8'hb3 == ex_bh_value ? pattern_table_179 : _GEN_690; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_692 = 8'hb4 == ex_bh_value ? pattern_table_180 : _GEN_691; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_693 = 8'hb5 == ex_bh_value ? pattern_table_181 : _GEN_692; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_694 = 8'hb6 == ex_bh_value ? pattern_table_182 : _GEN_693; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_695 = 8'hb7 == ex_bh_value ? pattern_table_183 : _GEN_694; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_696 = 8'hb8 == ex_bh_value ? pattern_table_184 : _GEN_695; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_697 = 8'hb9 == ex_bh_value ? pattern_table_185 : _GEN_696; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_698 = 8'hba == ex_bh_value ? pattern_table_186 : _GEN_697; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_699 = 8'hbb == ex_bh_value ? pattern_table_187 : _GEN_698; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_700 = 8'hbc == ex_bh_value ? pattern_table_188 : _GEN_699; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_701 = 8'hbd == ex_bh_value ? pattern_table_189 : _GEN_700; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_702 = 8'hbe == ex_bh_value ? pattern_table_190 : _GEN_701; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_703 = 8'hbf == ex_bh_value ? pattern_table_191 : _GEN_702; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_704 = 8'hc0 == ex_bh_value ? pattern_table_192 : _GEN_703; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_705 = 8'hc1 == ex_bh_value ? pattern_table_193 : _GEN_704; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_706 = 8'hc2 == ex_bh_value ? pattern_table_194 : _GEN_705; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_707 = 8'hc3 == ex_bh_value ? pattern_table_195 : _GEN_706; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_708 = 8'hc4 == ex_bh_value ? pattern_table_196 : _GEN_707; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_709 = 8'hc5 == ex_bh_value ? pattern_table_197 : _GEN_708; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_710 = 8'hc6 == ex_bh_value ? pattern_table_198 : _GEN_709; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_711 = 8'hc7 == ex_bh_value ? pattern_table_199 : _GEN_710; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_712 = 8'hc8 == ex_bh_value ? pattern_table_200 : _GEN_711; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_713 = 8'hc9 == ex_bh_value ? pattern_table_201 : _GEN_712; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_714 = 8'hca == ex_bh_value ? pattern_table_202 : _GEN_713; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_715 = 8'hcb == ex_bh_value ? pattern_table_203 : _GEN_714; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_716 = 8'hcc == ex_bh_value ? pattern_table_204 : _GEN_715; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_717 = 8'hcd == ex_bh_value ? pattern_table_205 : _GEN_716; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_718 = 8'hce == ex_bh_value ? pattern_table_206 : _GEN_717; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_719 = 8'hcf == ex_bh_value ? pattern_table_207 : _GEN_718; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_720 = 8'hd0 == ex_bh_value ? pattern_table_208 : _GEN_719; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_721 = 8'hd1 == ex_bh_value ? pattern_table_209 : _GEN_720; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_722 = 8'hd2 == ex_bh_value ? pattern_table_210 : _GEN_721; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_723 = 8'hd3 == ex_bh_value ? pattern_table_211 : _GEN_722; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_724 = 8'hd4 == ex_bh_value ? pattern_table_212 : _GEN_723; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_725 = 8'hd5 == ex_bh_value ? pattern_table_213 : _GEN_724; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_726 = 8'hd6 == ex_bh_value ? pattern_table_214 : _GEN_725; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_727 = 8'hd7 == ex_bh_value ? pattern_table_215 : _GEN_726; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_728 = 8'hd8 == ex_bh_value ? pattern_table_216 : _GEN_727; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_729 = 8'hd9 == ex_bh_value ? pattern_table_217 : _GEN_728; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_730 = 8'hda == ex_bh_value ? pattern_table_218 : _GEN_729; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_731 = 8'hdb == ex_bh_value ? pattern_table_219 : _GEN_730; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_732 = 8'hdc == ex_bh_value ? pattern_table_220 : _GEN_731; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_733 = 8'hdd == ex_bh_value ? pattern_table_221 : _GEN_732; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_734 = 8'hde == ex_bh_value ? pattern_table_222 : _GEN_733; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_735 = 8'hdf == ex_bh_value ? pattern_table_223 : _GEN_734; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_736 = 8'he0 == ex_bh_value ? pattern_table_224 : _GEN_735; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_737 = 8'he1 == ex_bh_value ? pattern_table_225 : _GEN_736; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_738 = 8'he2 == ex_bh_value ? pattern_table_226 : _GEN_737; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_739 = 8'he3 == ex_bh_value ? pattern_table_227 : _GEN_738; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_740 = 8'he4 == ex_bh_value ? pattern_table_228 : _GEN_739; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_741 = 8'he5 == ex_bh_value ? pattern_table_229 : _GEN_740; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_742 = 8'he6 == ex_bh_value ? pattern_table_230 : _GEN_741; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_743 = 8'he7 == ex_bh_value ? pattern_table_231 : _GEN_742; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_744 = 8'he8 == ex_bh_value ? pattern_table_232 : _GEN_743; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_745 = 8'he9 == ex_bh_value ? pattern_table_233 : _GEN_744; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_746 = 8'hea == ex_bh_value ? pattern_table_234 : _GEN_745; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_747 = 8'heb == ex_bh_value ? pattern_table_235 : _GEN_746; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_748 = 8'hec == ex_bh_value ? pattern_table_236 : _GEN_747; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_749 = 8'hed == ex_bh_value ? pattern_table_237 : _GEN_748; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_750 = 8'hee == ex_bh_value ? pattern_table_238 : _GEN_749; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_751 = 8'hef == ex_bh_value ? pattern_table_239 : _GEN_750; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_752 = 8'hf0 == ex_bh_value ? pattern_table_240 : _GEN_751; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_753 = 8'hf1 == ex_bh_value ? pattern_table_241 : _GEN_752; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_754 = 8'hf2 == ex_bh_value ? pattern_table_242 : _GEN_753; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_755 = 8'hf3 == ex_bh_value ? pattern_table_243 : _GEN_754; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_756 = 8'hf4 == ex_bh_value ? pattern_table_244 : _GEN_755; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_757 = 8'hf5 == ex_bh_value ? pattern_table_245 : _GEN_756; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_758 = 8'hf6 == ex_bh_value ? pattern_table_246 : _GEN_757; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_759 = 8'hf7 == ex_bh_value ? pattern_table_247 : _GEN_758; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_760 = 8'hf8 == ex_bh_value ? pattern_table_248 : _GEN_759; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_761 = 8'hf9 == ex_bh_value ? pattern_table_249 : _GEN_760; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_762 = 8'hfa == ex_bh_value ? pattern_table_250 : _GEN_761; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_763 = 8'hfb == ex_bh_value ? pattern_table_251 : _GEN_762; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_764 = 8'hfc == ex_bh_value ? pattern_table_252 : _GEN_763; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_765 = 8'hfd == ex_bh_value ? pattern_table_253 : _GEN_764; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_766 = 8'hfe == ex_bh_value ? pattern_table_254 : _GEN_765; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_767 = 8'hff == ex_bh_value ? pattern_table_255 : _GEN_766; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire  _pattern_table_T = 2'h0 == _GEN_767; // @[Conditional.scala 37:30]
  wire [1:0] _pattern_table_new_state_T = io_in_ex_io_br_io_br_flag ? 2'h1 : 2'h0; // @[BP.scala 79:39]
  wire  _pattern_table_T_1 = 2'h1 == _GEN_767; // @[Conditional.scala 37:30]
  wire [1:0] _pattern_table_new_state_T_1 = io_in_ex_io_br_io_br_flag ? 2'h2 : 2'h0; // @[BP.scala 80:39]
  wire  _pattern_table_T_2 = 2'h2 == _GEN_767; // @[Conditional.scala 37:30]
  wire [1:0] _pattern_table_new_state_T_2 = io_in_ex_io_br_io_br_flag ? 2'h3 : 2'h1; // @[BP.scala 81:39]
  wire  _pattern_table_T_3 = 2'h3 == _GEN_767; // @[Conditional.scala 37:30]
  wire [1:0] _pattern_table_new_state_T_3 = io_in_ex_io_br_io_br_flag ? 2'h3 : 2'h2; // @[BP.scala 82:39]
  wire [1:0] _GEN_768 = _pattern_table_T_3 ? _pattern_table_new_state_T_3 : 2'h1; // @[Conditional.scala 39:67 BP.scala 82:33]
  wire [1:0] _GEN_769 = _pattern_table_T_2 ? _pattern_table_new_state_T_2 : _GEN_768; // @[Conditional.scala 39:67 BP.scala 81:33]
  wire [1:0] _GEN_770 = _pattern_table_T_1 ? _pattern_table_new_state_T_1 : _GEN_769; // @[Conditional.scala 39:67 BP.scala 80:33]
  wire [7:0] bh_iodex = io_in_pc_io_reg_pc[9:2]; // @[BP.scala 100:29]
  wire [7:0] _GEN_2054 = 8'h1 == bh_iodex ? branch_history_1 : branch_history_0; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2055 = 8'h2 == bh_iodex ? branch_history_2 : _GEN_2054; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2056 = 8'h3 == bh_iodex ? branch_history_3 : _GEN_2055; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2057 = 8'h4 == bh_iodex ? branch_history_4 : _GEN_2056; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2058 = 8'h5 == bh_iodex ? branch_history_5 : _GEN_2057; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2059 = 8'h6 == bh_iodex ? branch_history_6 : _GEN_2058; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2060 = 8'h7 == bh_iodex ? branch_history_7 : _GEN_2059; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2061 = 8'h8 == bh_iodex ? branch_history_8 : _GEN_2060; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2062 = 8'h9 == bh_iodex ? branch_history_9 : _GEN_2061; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2063 = 8'ha == bh_iodex ? branch_history_10 : _GEN_2062; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2064 = 8'hb == bh_iodex ? branch_history_11 : _GEN_2063; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2065 = 8'hc == bh_iodex ? branch_history_12 : _GEN_2064; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2066 = 8'hd == bh_iodex ? branch_history_13 : _GEN_2065; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2067 = 8'he == bh_iodex ? branch_history_14 : _GEN_2066; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2068 = 8'hf == bh_iodex ? branch_history_15 : _GEN_2067; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2069 = 8'h10 == bh_iodex ? branch_history_16 : _GEN_2068; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2070 = 8'h11 == bh_iodex ? branch_history_17 : _GEN_2069; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2071 = 8'h12 == bh_iodex ? branch_history_18 : _GEN_2070; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2072 = 8'h13 == bh_iodex ? branch_history_19 : _GEN_2071; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2073 = 8'h14 == bh_iodex ? branch_history_20 : _GEN_2072; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2074 = 8'h15 == bh_iodex ? branch_history_21 : _GEN_2073; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2075 = 8'h16 == bh_iodex ? branch_history_22 : _GEN_2074; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2076 = 8'h17 == bh_iodex ? branch_history_23 : _GEN_2075; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2077 = 8'h18 == bh_iodex ? branch_history_24 : _GEN_2076; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2078 = 8'h19 == bh_iodex ? branch_history_25 : _GEN_2077; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2079 = 8'h1a == bh_iodex ? branch_history_26 : _GEN_2078; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2080 = 8'h1b == bh_iodex ? branch_history_27 : _GEN_2079; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2081 = 8'h1c == bh_iodex ? branch_history_28 : _GEN_2080; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2082 = 8'h1d == bh_iodex ? branch_history_29 : _GEN_2081; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2083 = 8'h1e == bh_iodex ? branch_history_30 : _GEN_2082; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2084 = 8'h1f == bh_iodex ? branch_history_31 : _GEN_2083; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2085 = 8'h20 == bh_iodex ? branch_history_32 : _GEN_2084; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2086 = 8'h21 == bh_iodex ? branch_history_33 : _GEN_2085; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2087 = 8'h22 == bh_iodex ? branch_history_34 : _GEN_2086; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2088 = 8'h23 == bh_iodex ? branch_history_35 : _GEN_2087; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2089 = 8'h24 == bh_iodex ? branch_history_36 : _GEN_2088; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2090 = 8'h25 == bh_iodex ? branch_history_37 : _GEN_2089; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2091 = 8'h26 == bh_iodex ? branch_history_38 : _GEN_2090; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2092 = 8'h27 == bh_iodex ? branch_history_39 : _GEN_2091; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2093 = 8'h28 == bh_iodex ? branch_history_40 : _GEN_2092; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2094 = 8'h29 == bh_iodex ? branch_history_41 : _GEN_2093; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2095 = 8'h2a == bh_iodex ? branch_history_42 : _GEN_2094; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2096 = 8'h2b == bh_iodex ? branch_history_43 : _GEN_2095; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2097 = 8'h2c == bh_iodex ? branch_history_44 : _GEN_2096; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2098 = 8'h2d == bh_iodex ? branch_history_45 : _GEN_2097; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2099 = 8'h2e == bh_iodex ? branch_history_46 : _GEN_2098; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2100 = 8'h2f == bh_iodex ? branch_history_47 : _GEN_2099; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2101 = 8'h30 == bh_iodex ? branch_history_48 : _GEN_2100; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2102 = 8'h31 == bh_iodex ? branch_history_49 : _GEN_2101; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2103 = 8'h32 == bh_iodex ? branch_history_50 : _GEN_2102; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2104 = 8'h33 == bh_iodex ? branch_history_51 : _GEN_2103; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2105 = 8'h34 == bh_iodex ? branch_history_52 : _GEN_2104; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2106 = 8'h35 == bh_iodex ? branch_history_53 : _GEN_2105; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2107 = 8'h36 == bh_iodex ? branch_history_54 : _GEN_2106; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2108 = 8'h37 == bh_iodex ? branch_history_55 : _GEN_2107; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2109 = 8'h38 == bh_iodex ? branch_history_56 : _GEN_2108; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2110 = 8'h39 == bh_iodex ? branch_history_57 : _GEN_2109; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2111 = 8'h3a == bh_iodex ? branch_history_58 : _GEN_2110; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2112 = 8'h3b == bh_iodex ? branch_history_59 : _GEN_2111; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2113 = 8'h3c == bh_iodex ? branch_history_60 : _GEN_2112; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2114 = 8'h3d == bh_iodex ? branch_history_61 : _GEN_2113; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2115 = 8'h3e == bh_iodex ? branch_history_62 : _GEN_2114; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2116 = 8'h3f == bh_iodex ? branch_history_63 : _GEN_2115; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2117 = 8'h40 == bh_iodex ? branch_history_64 : _GEN_2116; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2118 = 8'h41 == bh_iodex ? branch_history_65 : _GEN_2117; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2119 = 8'h42 == bh_iodex ? branch_history_66 : _GEN_2118; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2120 = 8'h43 == bh_iodex ? branch_history_67 : _GEN_2119; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2121 = 8'h44 == bh_iodex ? branch_history_68 : _GEN_2120; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2122 = 8'h45 == bh_iodex ? branch_history_69 : _GEN_2121; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2123 = 8'h46 == bh_iodex ? branch_history_70 : _GEN_2122; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2124 = 8'h47 == bh_iodex ? branch_history_71 : _GEN_2123; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2125 = 8'h48 == bh_iodex ? branch_history_72 : _GEN_2124; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2126 = 8'h49 == bh_iodex ? branch_history_73 : _GEN_2125; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2127 = 8'h4a == bh_iodex ? branch_history_74 : _GEN_2126; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2128 = 8'h4b == bh_iodex ? branch_history_75 : _GEN_2127; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2129 = 8'h4c == bh_iodex ? branch_history_76 : _GEN_2128; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2130 = 8'h4d == bh_iodex ? branch_history_77 : _GEN_2129; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2131 = 8'h4e == bh_iodex ? branch_history_78 : _GEN_2130; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2132 = 8'h4f == bh_iodex ? branch_history_79 : _GEN_2131; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2133 = 8'h50 == bh_iodex ? branch_history_80 : _GEN_2132; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2134 = 8'h51 == bh_iodex ? branch_history_81 : _GEN_2133; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2135 = 8'h52 == bh_iodex ? branch_history_82 : _GEN_2134; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2136 = 8'h53 == bh_iodex ? branch_history_83 : _GEN_2135; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2137 = 8'h54 == bh_iodex ? branch_history_84 : _GEN_2136; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2138 = 8'h55 == bh_iodex ? branch_history_85 : _GEN_2137; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2139 = 8'h56 == bh_iodex ? branch_history_86 : _GEN_2138; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2140 = 8'h57 == bh_iodex ? branch_history_87 : _GEN_2139; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2141 = 8'h58 == bh_iodex ? branch_history_88 : _GEN_2140; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2142 = 8'h59 == bh_iodex ? branch_history_89 : _GEN_2141; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2143 = 8'h5a == bh_iodex ? branch_history_90 : _GEN_2142; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2144 = 8'h5b == bh_iodex ? branch_history_91 : _GEN_2143; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2145 = 8'h5c == bh_iodex ? branch_history_92 : _GEN_2144; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2146 = 8'h5d == bh_iodex ? branch_history_93 : _GEN_2145; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2147 = 8'h5e == bh_iodex ? branch_history_94 : _GEN_2146; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2148 = 8'h5f == bh_iodex ? branch_history_95 : _GEN_2147; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2149 = 8'h60 == bh_iodex ? branch_history_96 : _GEN_2148; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2150 = 8'h61 == bh_iodex ? branch_history_97 : _GEN_2149; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2151 = 8'h62 == bh_iodex ? branch_history_98 : _GEN_2150; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2152 = 8'h63 == bh_iodex ? branch_history_99 : _GEN_2151; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2153 = 8'h64 == bh_iodex ? branch_history_100 : _GEN_2152; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2154 = 8'h65 == bh_iodex ? branch_history_101 : _GEN_2153; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2155 = 8'h66 == bh_iodex ? branch_history_102 : _GEN_2154; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2156 = 8'h67 == bh_iodex ? branch_history_103 : _GEN_2155; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2157 = 8'h68 == bh_iodex ? branch_history_104 : _GEN_2156; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2158 = 8'h69 == bh_iodex ? branch_history_105 : _GEN_2157; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2159 = 8'h6a == bh_iodex ? branch_history_106 : _GEN_2158; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2160 = 8'h6b == bh_iodex ? branch_history_107 : _GEN_2159; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2161 = 8'h6c == bh_iodex ? branch_history_108 : _GEN_2160; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2162 = 8'h6d == bh_iodex ? branch_history_109 : _GEN_2161; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2163 = 8'h6e == bh_iodex ? branch_history_110 : _GEN_2162; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2164 = 8'h6f == bh_iodex ? branch_history_111 : _GEN_2163; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2165 = 8'h70 == bh_iodex ? branch_history_112 : _GEN_2164; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2166 = 8'h71 == bh_iodex ? branch_history_113 : _GEN_2165; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2167 = 8'h72 == bh_iodex ? branch_history_114 : _GEN_2166; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2168 = 8'h73 == bh_iodex ? branch_history_115 : _GEN_2167; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2169 = 8'h74 == bh_iodex ? branch_history_116 : _GEN_2168; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2170 = 8'h75 == bh_iodex ? branch_history_117 : _GEN_2169; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2171 = 8'h76 == bh_iodex ? branch_history_118 : _GEN_2170; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2172 = 8'h77 == bh_iodex ? branch_history_119 : _GEN_2171; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2173 = 8'h78 == bh_iodex ? branch_history_120 : _GEN_2172; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2174 = 8'h79 == bh_iodex ? branch_history_121 : _GEN_2173; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2175 = 8'h7a == bh_iodex ? branch_history_122 : _GEN_2174; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2176 = 8'h7b == bh_iodex ? branch_history_123 : _GEN_2175; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2177 = 8'h7c == bh_iodex ? branch_history_124 : _GEN_2176; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2178 = 8'h7d == bh_iodex ? branch_history_125 : _GEN_2177; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2179 = 8'h7e == bh_iodex ? branch_history_126 : _GEN_2178; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2180 = 8'h7f == bh_iodex ? branch_history_127 : _GEN_2179; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2181 = 8'h80 == bh_iodex ? branch_history_128 : _GEN_2180; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2182 = 8'h81 == bh_iodex ? branch_history_129 : _GEN_2181; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2183 = 8'h82 == bh_iodex ? branch_history_130 : _GEN_2182; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2184 = 8'h83 == bh_iodex ? branch_history_131 : _GEN_2183; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2185 = 8'h84 == bh_iodex ? branch_history_132 : _GEN_2184; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2186 = 8'h85 == bh_iodex ? branch_history_133 : _GEN_2185; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2187 = 8'h86 == bh_iodex ? branch_history_134 : _GEN_2186; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2188 = 8'h87 == bh_iodex ? branch_history_135 : _GEN_2187; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2189 = 8'h88 == bh_iodex ? branch_history_136 : _GEN_2188; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2190 = 8'h89 == bh_iodex ? branch_history_137 : _GEN_2189; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2191 = 8'h8a == bh_iodex ? branch_history_138 : _GEN_2190; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2192 = 8'h8b == bh_iodex ? branch_history_139 : _GEN_2191; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2193 = 8'h8c == bh_iodex ? branch_history_140 : _GEN_2192; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2194 = 8'h8d == bh_iodex ? branch_history_141 : _GEN_2193; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2195 = 8'h8e == bh_iodex ? branch_history_142 : _GEN_2194; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2196 = 8'h8f == bh_iodex ? branch_history_143 : _GEN_2195; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2197 = 8'h90 == bh_iodex ? branch_history_144 : _GEN_2196; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2198 = 8'h91 == bh_iodex ? branch_history_145 : _GEN_2197; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2199 = 8'h92 == bh_iodex ? branch_history_146 : _GEN_2198; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2200 = 8'h93 == bh_iodex ? branch_history_147 : _GEN_2199; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2201 = 8'h94 == bh_iodex ? branch_history_148 : _GEN_2200; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2202 = 8'h95 == bh_iodex ? branch_history_149 : _GEN_2201; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2203 = 8'h96 == bh_iodex ? branch_history_150 : _GEN_2202; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2204 = 8'h97 == bh_iodex ? branch_history_151 : _GEN_2203; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2205 = 8'h98 == bh_iodex ? branch_history_152 : _GEN_2204; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2206 = 8'h99 == bh_iodex ? branch_history_153 : _GEN_2205; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2207 = 8'h9a == bh_iodex ? branch_history_154 : _GEN_2206; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2208 = 8'h9b == bh_iodex ? branch_history_155 : _GEN_2207; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2209 = 8'h9c == bh_iodex ? branch_history_156 : _GEN_2208; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2210 = 8'h9d == bh_iodex ? branch_history_157 : _GEN_2209; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2211 = 8'h9e == bh_iodex ? branch_history_158 : _GEN_2210; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2212 = 8'h9f == bh_iodex ? branch_history_159 : _GEN_2211; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2213 = 8'ha0 == bh_iodex ? branch_history_160 : _GEN_2212; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2214 = 8'ha1 == bh_iodex ? branch_history_161 : _GEN_2213; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2215 = 8'ha2 == bh_iodex ? branch_history_162 : _GEN_2214; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2216 = 8'ha3 == bh_iodex ? branch_history_163 : _GEN_2215; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2217 = 8'ha4 == bh_iodex ? branch_history_164 : _GEN_2216; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2218 = 8'ha5 == bh_iodex ? branch_history_165 : _GEN_2217; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2219 = 8'ha6 == bh_iodex ? branch_history_166 : _GEN_2218; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2220 = 8'ha7 == bh_iodex ? branch_history_167 : _GEN_2219; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2221 = 8'ha8 == bh_iodex ? branch_history_168 : _GEN_2220; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2222 = 8'ha9 == bh_iodex ? branch_history_169 : _GEN_2221; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2223 = 8'haa == bh_iodex ? branch_history_170 : _GEN_2222; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2224 = 8'hab == bh_iodex ? branch_history_171 : _GEN_2223; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2225 = 8'hac == bh_iodex ? branch_history_172 : _GEN_2224; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2226 = 8'had == bh_iodex ? branch_history_173 : _GEN_2225; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2227 = 8'hae == bh_iodex ? branch_history_174 : _GEN_2226; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2228 = 8'haf == bh_iodex ? branch_history_175 : _GEN_2227; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2229 = 8'hb0 == bh_iodex ? branch_history_176 : _GEN_2228; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2230 = 8'hb1 == bh_iodex ? branch_history_177 : _GEN_2229; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2231 = 8'hb2 == bh_iodex ? branch_history_178 : _GEN_2230; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2232 = 8'hb3 == bh_iodex ? branch_history_179 : _GEN_2231; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2233 = 8'hb4 == bh_iodex ? branch_history_180 : _GEN_2232; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2234 = 8'hb5 == bh_iodex ? branch_history_181 : _GEN_2233; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2235 = 8'hb6 == bh_iodex ? branch_history_182 : _GEN_2234; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2236 = 8'hb7 == bh_iodex ? branch_history_183 : _GEN_2235; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2237 = 8'hb8 == bh_iodex ? branch_history_184 : _GEN_2236; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2238 = 8'hb9 == bh_iodex ? branch_history_185 : _GEN_2237; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2239 = 8'hba == bh_iodex ? branch_history_186 : _GEN_2238; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2240 = 8'hbb == bh_iodex ? branch_history_187 : _GEN_2239; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2241 = 8'hbc == bh_iodex ? branch_history_188 : _GEN_2240; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2242 = 8'hbd == bh_iodex ? branch_history_189 : _GEN_2241; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2243 = 8'hbe == bh_iodex ? branch_history_190 : _GEN_2242; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2244 = 8'hbf == bh_iodex ? branch_history_191 : _GEN_2243; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2245 = 8'hc0 == bh_iodex ? branch_history_192 : _GEN_2244; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2246 = 8'hc1 == bh_iodex ? branch_history_193 : _GEN_2245; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2247 = 8'hc2 == bh_iodex ? branch_history_194 : _GEN_2246; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2248 = 8'hc3 == bh_iodex ? branch_history_195 : _GEN_2247; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2249 = 8'hc4 == bh_iodex ? branch_history_196 : _GEN_2248; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2250 = 8'hc5 == bh_iodex ? branch_history_197 : _GEN_2249; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2251 = 8'hc6 == bh_iodex ? branch_history_198 : _GEN_2250; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2252 = 8'hc7 == bh_iodex ? branch_history_199 : _GEN_2251; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2253 = 8'hc8 == bh_iodex ? branch_history_200 : _GEN_2252; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2254 = 8'hc9 == bh_iodex ? branch_history_201 : _GEN_2253; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2255 = 8'hca == bh_iodex ? branch_history_202 : _GEN_2254; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2256 = 8'hcb == bh_iodex ? branch_history_203 : _GEN_2255; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2257 = 8'hcc == bh_iodex ? branch_history_204 : _GEN_2256; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2258 = 8'hcd == bh_iodex ? branch_history_205 : _GEN_2257; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2259 = 8'hce == bh_iodex ? branch_history_206 : _GEN_2258; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2260 = 8'hcf == bh_iodex ? branch_history_207 : _GEN_2259; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2261 = 8'hd0 == bh_iodex ? branch_history_208 : _GEN_2260; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2262 = 8'hd1 == bh_iodex ? branch_history_209 : _GEN_2261; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2263 = 8'hd2 == bh_iodex ? branch_history_210 : _GEN_2262; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2264 = 8'hd3 == bh_iodex ? branch_history_211 : _GEN_2263; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2265 = 8'hd4 == bh_iodex ? branch_history_212 : _GEN_2264; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2266 = 8'hd5 == bh_iodex ? branch_history_213 : _GEN_2265; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2267 = 8'hd6 == bh_iodex ? branch_history_214 : _GEN_2266; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2268 = 8'hd7 == bh_iodex ? branch_history_215 : _GEN_2267; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2269 = 8'hd8 == bh_iodex ? branch_history_216 : _GEN_2268; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2270 = 8'hd9 == bh_iodex ? branch_history_217 : _GEN_2269; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2271 = 8'hda == bh_iodex ? branch_history_218 : _GEN_2270; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2272 = 8'hdb == bh_iodex ? branch_history_219 : _GEN_2271; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2273 = 8'hdc == bh_iodex ? branch_history_220 : _GEN_2272; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2274 = 8'hdd == bh_iodex ? branch_history_221 : _GEN_2273; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2275 = 8'hde == bh_iodex ? branch_history_222 : _GEN_2274; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2276 = 8'hdf == bh_iodex ? branch_history_223 : _GEN_2275; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2277 = 8'he0 == bh_iodex ? branch_history_224 : _GEN_2276; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2278 = 8'he1 == bh_iodex ? branch_history_225 : _GEN_2277; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2279 = 8'he2 == bh_iodex ? branch_history_226 : _GEN_2278; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2280 = 8'he3 == bh_iodex ? branch_history_227 : _GEN_2279; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2281 = 8'he4 == bh_iodex ? branch_history_228 : _GEN_2280; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2282 = 8'he5 == bh_iodex ? branch_history_229 : _GEN_2281; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2283 = 8'he6 == bh_iodex ? branch_history_230 : _GEN_2282; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2284 = 8'he7 == bh_iodex ? branch_history_231 : _GEN_2283; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2285 = 8'he8 == bh_iodex ? branch_history_232 : _GEN_2284; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2286 = 8'he9 == bh_iodex ? branch_history_233 : _GEN_2285; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2287 = 8'hea == bh_iodex ? branch_history_234 : _GEN_2286; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2288 = 8'heb == bh_iodex ? branch_history_235 : _GEN_2287; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2289 = 8'hec == bh_iodex ? branch_history_236 : _GEN_2288; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2290 = 8'hed == bh_iodex ? branch_history_237 : _GEN_2289; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2291 = 8'hee == bh_iodex ? branch_history_238 : _GEN_2290; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2292 = 8'hef == bh_iodex ? branch_history_239 : _GEN_2291; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2293 = 8'hf0 == bh_iodex ? branch_history_240 : _GEN_2292; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2294 = 8'hf1 == bh_iodex ? branch_history_241 : _GEN_2293; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2295 = 8'hf2 == bh_iodex ? branch_history_242 : _GEN_2294; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2296 = 8'hf3 == bh_iodex ? branch_history_243 : _GEN_2295; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2297 = 8'hf4 == bh_iodex ? branch_history_244 : _GEN_2296; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2298 = 8'hf5 == bh_iodex ? branch_history_245 : _GEN_2297; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2299 = 8'hf6 == bh_iodex ? branch_history_246 : _GEN_2298; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2300 = 8'hf7 == bh_iodex ? branch_history_247 : _GEN_2299; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2301 = 8'hf8 == bh_iodex ? branch_history_248 : _GEN_2300; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2302 = 8'hf9 == bh_iodex ? branch_history_249 : _GEN_2301; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2303 = 8'hfa == bh_iodex ? branch_history_250 : _GEN_2302; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2304 = 8'hfb == bh_iodex ? branch_history_251 : _GEN_2303; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2305 = 8'hfc == bh_iodex ? branch_history_252 : _GEN_2304; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2306 = 8'hfd == bh_iodex ? branch_history_253 : _GEN_2305; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] _GEN_2307 = 8'hfe == bh_iodex ? branch_history_254 : _GEN_2306; // @[BP.scala 101:48 BP.scala 101:48]
  wire [7:0] bh_value = 8'hff == bh_iodex ? branch_history_255 : _GEN_2307; // @[BP.scala 101:48 BP.scala 101:48]
  wire [31:0] _pt_flag_T = io_in_pc_io_inst & 32'h707f; // @[BP.scala 107:15]
  wire  _pt_flag_T_1 = 32'h63 == _pt_flag_T; // @[BP.scala 107:15]
  wire  _pt_flag_T_3 = 32'h1063 == _pt_flag_T; // @[BP.scala 108:15]
  wire  _pt_flag_T_5 = 32'h5063 == _pt_flag_T; // @[BP.scala 109:15]
  wire  _pt_flag_T_7 = 32'h7063 == _pt_flag_T; // @[BP.scala 110:15]
  wire  _pt_flag_T_9 = 32'h4063 == _pt_flag_T; // @[BP.scala 111:15]
  wire  _pt_flag_T_11 = 32'h6063 == _pt_flag_T; // @[BP.scala 112:15]
  wire  pt_flag = _pt_flag_T_1 | (_pt_flag_T_3 | (_pt_flag_T_5 | (_pt_flag_T_7 | (_pt_flag_T_9 | _pt_flag_T_11)))); // @[Mux.scala 98:16]
  wire [1:0] _GEN_2310 = 8'h1 == bh_value ? pattern_table_1 : pattern_table_0; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2311 = 8'h2 == bh_value ? pattern_table_2 : _GEN_2310; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2312 = 8'h3 == bh_value ? pattern_table_3 : _GEN_2311; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2313 = 8'h4 == bh_value ? pattern_table_4 : _GEN_2312; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2314 = 8'h5 == bh_value ? pattern_table_5 : _GEN_2313; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2315 = 8'h6 == bh_value ? pattern_table_6 : _GEN_2314; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2316 = 8'h7 == bh_value ? pattern_table_7 : _GEN_2315; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2317 = 8'h8 == bh_value ? pattern_table_8 : _GEN_2316; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2318 = 8'h9 == bh_value ? pattern_table_9 : _GEN_2317; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2319 = 8'ha == bh_value ? pattern_table_10 : _GEN_2318; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2320 = 8'hb == bh_value ? pattern_table_11 : _GEN_2319; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2321 = 8'hc == bh_value ? pattern_table_12 : _GEN_2320; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2322 = 8'hd == bh_value ? pattern_table_13 : _GEN_2321; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2323 = 8'he == bh_value ? pattern_table_14 : _GEN_2322; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2324 = 8'hf == bh_value ? pattern_table_15 : _GEN_2323; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2325 = 8'h10 == bh_value ? pattern_table_16 : _GEN_2324; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2326 = 8'h11 == bh_value ? pattern_table_17 : _GEN_2325; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2327 = 8'h12 == bh_value ? pattern_table_18 : _GEN_2326; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2328 = 8'h13 == bh_value ? pattern_table_19 : _GEN_2327; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2329 = 8'h14 == bh_value ? pattern_table_20 : _GEN_2328; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2330 = 8'h15 == bh_value ? pattern_table_21 : _GEN_2329; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2331 = 8'h16 == bh_value ? pattern_table_22 : _GEN_2330; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2332 = 8'h17 == bh_value ? pattern_table_23 : _GEN_2331; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2333 = 8'h18 == bh_value ? pattern_table_24 : _GEN_2332; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2334 = 8'h19 == bh_value ? pattern_table_25 : _GEN_2333; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2335 = 8'h1a == bh_value ? pattern_table_26 : _GEN_2334; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2336 = 8'h1b == bh_value ? pattern_table_27 : _GEN_2335; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2337 = 8'h1c == bh_value ? pattern_table_28 : _GEN_2336; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2338 = 8'h1d == bh_value ? pattern_table_29 : _GEN_2337; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2339 = 8'h1e == bh_value ? pattern_table_30 : _GEN_2338; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2340 = 8'h1f == bh_value ? pattern_table_31 : _GEN_2339; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2341 = 8'h20 == bh_value ? pattern_table_32 : _GEN_2340; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2342 = 8'h21 == bh_value ? pattern_table_33 : _GEN_2341; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2343 = 8'h22 == bh_value ? pattern_table_34 : _GEN_2342; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2344 = 8'h23 == bh_value ? pattern_table_35 : _GEN_2343; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2345 = 8'h24 == bh_value ? pattern_table_36 : _GEN_2344; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2346 = 8'h25 == bh_value ? pattern_table_37 : _GEN_2345; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2347 = 8'h26 == bh_value ? pattern_table_38 : _GEN_2346; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2348 = 8'h27 == bh_value ? pattern_table_39 : _GEN_2347; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2349 = 8'h28 == bh_value ? pattern_table_40 : _GEN_2348; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2350 = 8'h29 == bh_value ? pattern_table_41 : _GEN_2349; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2351 = 8'h2a == bh_value ? pattern_table_42 : _GEN_2350; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2352 = 8'h2b == bh_value ? pattern_table_43 : _GEN_2351; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2353 = 8'h2c == bh_value ? pattern_table_44 : _GEN_2352; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2354 = 8'h2d == bh_value ? pattern_table_45 : _GEN_2353; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2355 = 8'h2e == bh_value ? pattern_table_46 : _GEN_2354; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2356 = 8'h2f == bh_value ? pattern_table_47 : _GEN_2355; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2357 = 8'h30 == bh_value ? pattern_table_48 : _GEN_2356; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2358 = 8'h31 == bh_value ? pattern_table_49 : _GEN_2357; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2359 = 8'h32 == bh_value ? pattern_table_50 : _GEN_2358; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2360 = 8'h33 == bh_value ? pattern_table_51 : _GEN_2359; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2361 = 8'h34 == bh_value ? pattern_table_52 : _GEN_2360; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2362 = 8'h35 == bh_value ? pattern_table_53 : _GEN_2361; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2363 = 8'h36 == bh_value ? pattern_table_54 : _GEN_2362; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2364 = 8'h37 == bh_value ? pattern_table_55 : _GEN_2363; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2365 = 8'h38 == bh_value ? pattern_table_56 : _GEN_2364; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2366 = 8'h39 == bh_value ? pattern_table_57 : _GEN_2365; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2367 = 8'h3a == bh_value ? pattern_table_58 : _GEN_2366; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2368 = 8'h3b == bh_value ? pattern_table_59 : _GEN_2367; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2369 = 8'h3c == bh_value ? pattern_table_60 : _GEN_2368; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2370 = 8'h3d == bh_value ? pattern_table_61 : _GEN_2369; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2371 = 8'h3e == bh_value ? pattern_table_62 : _GEN_2370; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2372 = 8'h3f == bh_value ? pattern_table_63 : _GEN_2371; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2373 = 8'h40 == bh_value ? pattern_table_64 : _GEN_2372; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2374 = 8'h41 == bh_value ? pattern_table_65 : _GEN_2373; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2375 = 8'h42 == bh_value ? pattern_table_66 : _GEN_2374; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2376 = 8'h43 == bh_value ? pattern_table_67 : _GEN_2375; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2377 = 8'h44 == bh_value ? pattern_table_68 : _GEN_2376; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2378 = 8'h45 == bh_value ? pattern_table_69 : _GEN_2377; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2379 = 8'h46 == bh_value ? pattern_table_70 : _GEN_2378; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2380 = 8'h47 == bh_value ? pattern_table_71 : _GEN_2379; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2381 = 8'h48 == bh_value ? pattern_table_72 : _GEN_2380; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2382 = 8'h49 == bh_value ? pattern_table_73 : _GEN_2381; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2383 = 8'h4a == bh_value ? pattern_table_74 : _GEN_2382; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2384 = 8'h4b == bh_value ? pattern_table_75 : _GEN_2383; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2385 = 8'h4c == bh_value ? pattern_table_76 : _GEN_2384; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2386 = 8'h4d == bh_value ? pattern_table_77 : _GEN_2385; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2387 = 8'h4e == bh_value ? pattern_table_78 : _GEN_2386; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2388 = 8'h4f == bh_value ? pattern_table_79 : _GEN_2387; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2389 = 8'h50 == bh_value ? pattern_table_80 : _GEN_2388; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2390 = 8'h51 == bh_value ? pattern_table_81 : _GEN_2389; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2391 = 8'h52 == bh_value ? pattern_table_82 : _GEN_2390; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2392 = 8'h53 == bh_value ? pattern_table_83 : _GEN_2391; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2393 = 8'h54 == bh_value ? pattern_table_84 : _GEN_2392; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2394 = 8'h55 == bh_value ? pattern_table_85 : _GEN_2393; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2395 = 8'h56 == bh_value ? pattern_table_86 : _GEN_2394; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2396 = 8'h57 == bh_value ? pattern_table_87 : _GEN_2395; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2397 = 8'h58 == bh_value ? pattern_table_88 : _GEN_2396; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2398 = 8'h59 == bh_value ? pattern_table_89 : _GEN_2397; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2399 = 8'h5a == bh_value ? pattern_table_90 : _GEN_2398; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2400 = 8'h5b == bh_value ? pattern_table_91 : _GEN_2399; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2401 = 8'h5c == bh_value ? pattern_table_92 : _GEN_2400; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2402 = 8'h5d == bh_value ? pattern_table_93 : _GEN_2401; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2403 = 8'h5e == bh_value ? pattern_table_94 : _GEN_2402; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2404 = 8'h5f == bh_value ? pattern_table_95 : _GEN_2403; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2405 = 8'h60 == bh_value ? pattern_table_96 : _GEN_2404; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2406 = 8'h61 == bh_value ? pattern_table_97 : _GEN_2405; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2407 = 8'h62 == bh_value ? pattern_table_98 : _GEN_2406; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2408 = 8'h63 == bh_value ? pattern_table_99 : _GEN_2407; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2409 = 8'h64 == bh_value ? pattern_table_100 : _GEN_2408; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2410 = 8'h65 == bh_value ? pattern_table_101 : _GEN_2409; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2411 = 8'h66 == bh_value ? pattern_table_102 : _GEN_2410; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2412 = 8'h67 == bh_value ? pattern_table_103 : _GEN_2411; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2413 = 8'h68 == bh_value ? pattern_table_104 : _GEN_2412; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2414 = 8'h69 == bh_value ? pattern_table_105 : _GEN_2413; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2415 = 8'h6a == bh_value ? pattern_table_106 : _GEN_2414; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2416 = 8'h6b == bh_value ? pattern_table_107 : _GEN_2415; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2417 = 8'h6c == bh_value ? pattern_table_108 : _GEN_2416; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2418 = 8'h6d == bh_value ? pattern_table_109 : _GEN_2417; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2419 = 8'h6e == bh_value ? pattern_table_110 : _GEN_2418; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2420 = 8'h6f == bh_value ? pattern_table_111 : _GEN_2419; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2421 = 8'h70 == bh_value ? pattern_table_112 : _GEN_2420; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2422 = 8'h71 == bh_value ? pattern_table_113 : _GEN_2421; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2423 = 8'h72 == bh_value ? pattern_table_114 : _GEN_2422; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2424 = 8'h73 == bh_value ? pattern_table_115 : _GEN_2423; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2425 = 8'h74 == bh_value ? pattern_table_116 : _GEN_2424; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2426 = 8'h75 == bh_value ? pattern_table_117 : _GEN_2425; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2427 = 8'h76 == bh_value ? pattern_table_118 : _GEN_2426; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2428 = 8'h77 == bh_value ? pattern_table_119 : _GEN_2427; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2429 = 8'h78 == bh_value ? pattern_table_120 : _GEN_2428; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2430 = 8'h79 == bh_value ? pattern_table_121 : _GEN_2429; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2431 = 8'h7a == bh_value ? pattern_table_122 : _GEN_2430; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2432 = 8'h7b == bh_value ? pattern_table_123 : _GEN_2431; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2433 = 8'h7c == bh_value ? pattern_table_124 : _GEN_2432; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2434 = 8'h7d == bh_value ? pattern_table_125 : _GEN_2433; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2435 = 8'h7e == bh_value ? pattern_table_126 : _GEN_2434; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2436 = 8'h7f == bh_value ? pattern_table_127 : _GEN_2435; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2437 = 8'h80 == bh_value ? pattern_table_128 : _GEN_2436; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2438 = 8'h81 == bh_value ? pattern_table_129 : _GEN_2437; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2439 = 8'h82 == bh_value ? pattern_table_130 : _GEN_2438; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2440 = 8'h83 == bh_value ? pattern_table_131 : _GEN_2439; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2441 = 8'h84 == bh_value ? pattern_table_132 : _GEN_2440; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2442 = 8'h85 == bh_value ? pattern_table_133 : _GEN_2441; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2443 = 8'h86 == bh_value ? pattern_table_134 : _GEN_2442; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2444 = 8'h87 == bh_value ? pattern_table_135 : _GEN_2443; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2445 = 8'h88 == bh_value ? pattern_table_136 : _GEN_2444; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2446 = 8'h89 == bh_value ? pattern_table_137 : _GEN_2445; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2447 = 8'h8a == bh_value ? pattern_table_138 : _GEN_2446; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2448 = 8'h8b == bh_value ? pattern_table_139 : _GEN_2447; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2449 = 8'h8c == bh_value ? pattern_table_140 : _GEN_2448; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2450 = 8'h8d == bh_value ? pattern_table_141 : _GEN_2449; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2451 = 8'h8e == bh_value ? pattern_table_142 : _GEN_2450; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2452 = 8'h8f == bh_value ? pattern_table_143 : _GEN_2451; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2453 = 8'h90 == bh_value ? pattern_table_144 : _GEN_2452; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2454 = 8'h91 == bh_value ? pattern_table_145 : _GEN_2453; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2455 = 8'h92 == bh_value ? pattern_table_146 : _GEN_2454; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2456 = 8'h93 == bh_value ? pattern_table_147 : _GEN_2455; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2457 = 8'h94 == bh_value ? pattern_table_148 : _GEN_2456; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2458 = 8'h95 == bh_value ? pattern_table_149 : _GEN_2457; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2459 = 8'h96 == bh_value ? pattern_table_150 : _GEN_2458; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2460 = 8'h97 == bh_value ? pattern_table_151 : _GEN_2459; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2461 = 8'h98 == bh_value ? pattern_table_152 : _GEN_2460; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2462 = 8'h99 == bh_value ? pattern_table_153 : _GEN_2461; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2463 = 8'h9a == bh_value ? pattern_table_154 : _GEN_2462; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2464 = 8'h9b == bh_value ? pattern_table_155 : _GEN_2463; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2465 = 8'h9c == bh_value ? pattern_table_156 : _GEN_2464; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2466 = 8'h9d == bh_value ? pattern_table_157 : _GEN_2465; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2467 = 8'h9e == bh_value ? pattern_table_158 : _GEN_2466; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2468 = 8'h9f == bh_value ? pattern_table_159 : _GEN_2467; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2469 = 8'ha0 == bh_value ? pattern_table_160 : _GEN_2468; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2470 = 8'ha1 == bh_value ? pattern_table_161 : _GEN_2469; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2471 = 8'ha2 == bh_value ? pattern_table_162 : _GEN_2470; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2472 = 8'ha3 == bh_value ? pattern_table_163 : _GEN_2471; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2473 = 8'ha4 == bh_value ? pattern_table_164 : _GEN_2472; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2474 = 8'ha5 == bh_value ? pattern_table_165 : _GEN_2473; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2475 = 8'ha6 == bh_value ? pattern_table_166 : _GEN_2474; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2476 = 8'ha7 == bh_value ? pattern_table_167 : _GEN_2475; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2477 = 8'ha8 == bh_value ? pattern_table_168 : _GEN_2476; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2478 = 8'ha9 == bh_value ? pattern_table_169 : _GEN_2477; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2479 = 8'haa == bh_value ? pattern_table_170 : _GEN_2478; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2480 = 8'hab == bh_value ? pattern_table_171 : _GEN_2479; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2481 = 8'hac == bh_value ? pattern_table_172 : _GEN_2480; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2482 = 8'had == bh_value ? pattern_table_173 : _GEN_2481; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2483 = 8'hae == bh_value ? pattern_table_174 : _GEN_2482; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2484 = 8'haf == bh_value ? pattern_table_175 : _GEN_2483; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2485 = 8'hb0 == bh_value ? pattern_table_176 : _GEN_2484; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2486 = 8'hb1 == bh_value ? pattern_table_177 : _GEN_2485; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2487 = 8'hb2 == bh_value ? pattern_table_178 : _GEN_2486; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2488 = 8'hb3 == bh_value ? pattern_table_179 : _GEN_2487; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2489 = 8'hb4 == bh_value ? pattern_table_180 : _GEN_2488; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2490 = 8'hb5 == bh_value ? pattern_table_181 : _GEN_2489; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2491 = 8'hb6 == bh_value ? pattern_table_182 : _GEN_2490; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2492 = 8'hb7 == bh_value ? pattern_table_183 : _GEN_2491; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2493 = 8'hb8 == bh_value ? pattern_table_184 : _GEN_2492; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2494 = 8'hb9 == bh_value ? pattern_table_185 : _GEN_2493; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2495 = 8'hba == bh_value ? pattern_table_186 : _GEN_2494; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2496 = 8'hbb == bh_value ? pattern_table_187 : _GEN_2495; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2497 = 8'hbc == bh_value ? pattern_table_188 : _GEN_2496; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2498 = 8'hbd == bh_value ? pattern_table_189 : _GEN_2497; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2499 = 8'hbe == bh_value ? pattern_table_190 : _GEN_2498; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2500 = 8'hbf == bh_value ? pattern_table_191 : _GEN_2499; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2501 = 8'hc0 == bh_value ? pattern_table_192 : _GEN_2500; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2502 = 8'hc1 == bh_value ? pattern_table_193 : _GEN_2501; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2503 = 8'hc2 == bh_value ? pattern_table_194 : _GEN_2502; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2504 = 8'hc3 == bh_value ? pattern_table_195 : _GEN_2503; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2505 = 8'hc4 == bh_value ? pattern_table_196 : _GEN_2504; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2506 = 8'hc5 == bh_value ? pattern_table_197 : _GEN_2505; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2507 = 8'hc6 == bh_value ? pattern_table_198 : _GEN_2506; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2508 = 8'hc7 == bh_value ? pattern_table_199 : _GEN_2507; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2509 = 8'hc8 == bh_value ? pattern_table_200 : _GEN_2508; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2510 = 8'hc9 == bh_value ? pattern_table_201 : _GEN_2509; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2511 = 8'hca == bh_value ? pattern_table_202 : _GEN_2510; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2512 = 8'hcb == bh_value ? pattern_table_203 : _GEN_2511; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2513 = 8'hcc == bh_value ? pattern_table_204 : _GEN_2512; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2514 = 8'hcd == bh_value ? pattern_table_205 : _GEN_2513; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2515 = 8'hce == bh_value ? pattern_table_206 : _GEN_2514; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2516 = 8'hcf == bh_value ? pattern_table_207 : _GEN_2515; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2517 = 8'hd0 == bh_value ? pattern_table_208 : _GEN_2516; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2518 = 8'hd1 == bh_value ? pattern_table_209 : _GEN_2517; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2519 = 8'hd2 == bh_value ? pattern_table_210 : _GEN_2518; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2520 = 8'hd3 == bh_value ? pattern_table_211 : _GEN_2519; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2521 = 8'hd4 == bh_value ? pattern_table_212 : _GEN_2520; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2522 = 8'hd5 == bh_value ? pattern_table_213 : _GEN_2521; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2523 = 8'hd6 == bh_value ? pattern_table_214 : _GEN_2522; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2524 = 8'hd7 == bh_value ? pattern_table_215 : _GEN_2523; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2525 = 8'hd8 == bh_value ? pattern_table_216 : _GEN_2524; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2526 = 8'hd9 == bh_value ? pattern_table_217 : _GEN_2525; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2527 = 8'hda == bh_value ? pattern_table_218 : _GEN_2526; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2528 = 8'hdb == bh_value ? pattern_table_219 : _GEN_2527; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2529 = 8'hdc == bh_value ? pattern_table_220 : _GEN_2528; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2530 = 8'hdd == bh_value ? pattern_table_221 : _GEN_2529; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2531 = 8'hde == bh_value ? pattern_table_222 : _GEN_2530; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2532 = 8'hdf == bh_value ? pattern_table_223 : _GEN_2531; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2533 = 8'he0 == bh_value ? pattern_table_224 : _GEN_2532; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2534 = 8'he1 == bh_value ? pattern_table_225 : _GEN_2533; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2535 = 8'he2 == bh_value ? pattern_table_226 : _GEN_2534; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2536 = 8'he3 == bh_value ? pattern_table_227 : _GEN_2535; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2537 = 8'he4 == bh_value ? pattern_table_228 : _GEN_2536; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2538 = 8'he5 == bh_value ? pattern_table_229 : _GEN_2537; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2539 = 8'he6 == bh_value ? pattern_table_230 : _GEN_2538; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2540 = 8'he7 == bh_value ? pattern_table_231 : _GEN_2539; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2541 = 8'he8 == bh_value ? pattern_table_232 : _GEN_2540; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2542 = 8'he9 == bh_value ? pattern_table_233 : _GEN_2541; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2543 = 8'hea == bh_value ? pattern_table_234 : _GEN_2542; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2544 = 8'heb == bh_value ? pattern_table_235 : _GEN_2543; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2545 = 8'hec == bh_value ? pattern_table_236 : _GEN_2544; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2546 = 8'hed == bh_value ? pattern_table_237 : _GEN_2545; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2547 = 8'hee == bh_value ? pattern_table_238 : _GEN_2546; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2548 = 8'hef == bh_value ? pattern_table_239 : _GEN_2547; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2549 = 8'hf0 == bh_value ? pattern_table_240 : _GEN_2548; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2550 = 8'hf1 == bh_value ? pattern_table_241 : _GEN_2549; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2551 = 8'hf2 == bh_value ? pattern_table_242 : _GEN_2550; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2552 = 8'hf3 == bh_value ? pattern_table_243 : _GEN_2551; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2553 = 8'hf4 == bh_value ? pattern_table_244 : _GEN_2552; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2554 = 8'hf5 == bh_value ? pattern_table_245 : _GEN_2553; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2555 = 8'hf6 == bh_value ? pattern_table_246 : _GEN_2554; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2556 = 8'hf7 == bh_value ? pattern_table_247 : _GEN_2555; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2557 = 8'hf8 == bh_value ? pattern_table_248 : _GEN_2556; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2558 = 8'hf9 == bh_value ? pattern_table_249 : _GEN_2557; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2559 = 8'hfa == bh_value ? pattern_table_250 : _GEN_2558; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2560 = 8'hfb == bh_value ? pattern_table_251 : _GEN_2559; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2561 = 8'hfc == bh_value ? pattern_table_252 : _GEN_2560; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2562 = 8'hfd == bh_value ? pattern_table_253 : _GEN_2561; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2563 = 8'hfe == bh_value ? pattern_table_254 : _GEN_2562; // @[BP.scala 115:23 BP.scala 115:23]
  wire [1:0] _GEN_2564 = 8'hff == bh_value ? pattern_table_255 : _GEN_2563; // @[BP.scala 115:23 BP.scala 115:23]
  wire  _T_5 = _GEN_2564 == 2'h2 | _GEN_2564 == 2'h3; // @[BP.scala 115:30]
  wire [31:0] _T_6 = io_in_pc_io_inst & 32'h7f; // @[BP.scala 121:19]
  wire  _T_10 = 32'h6f == _T_6 | 32'h67 == _pt_flag_T; // @[BP.scala 121:27]
  wire  pred_flag = pt_flag ? _T_5 : _T_10; // @[BP.scala 114:19]
  wire [31:0] _GEN_2569 = 8'h1 == bh_iodex ? branch_target_buffer_1 : branch_target_buffer_0; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2570 = 8'h2 == bh_iodex ? branch_target_buffer_2 : _GEN_2569; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2571 = 8'h3 == bh_iodex ? branch_target_buffer_3 : _GEN_2570; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2572 = 8'h4 == bh_iodex ? branch_target_buffer_4 : _GEN_2571; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2573 = 8'h5 == bh_iodex ? branch_target_buffer_5 : _GEN_2572; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2574 = 8'h6 == bh_iodex ? branch_target_buffer_6 : _GEN_2573; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2575 = 8'h7 == bh_iodex ? branch_target_buffer_7 : _GEN_2574; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2576 = 8'h8 == bh_iodex ? branch_target_buffer_8 : _GEN_2575; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2577 = 8'h9 == bh_iodex ? branch_target_buffer_9 : _GEN_2576; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2578 = 8'ha == bh_iodex ? branch_target_buffer_10 : _GEN_2577; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2579 = 8'hb == bh_iodex ? branch_target_buffer_11 : _GEN_2578; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2580 = 8'hc == bh_iodex ? branch_target_buffer_12 : _GEN_2579; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2581 = 8'hd == bh_iodex ? branch_target_buffer_13 : _GEN_2580; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2582 = 8'he == bh_iodex ? branch_target_buffer_14 : _GEN_2581; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2583 = 8'hf == bh_iodex ? branch_target_buffer_15 : _GEN_2582; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2584 = 8'h10 == bh_iodex ? branch_target_buffer_16 : _GEN_2583; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2585 = 8'h11 == bh_iodex ? branch_target_buffer_17 : _GEN_2584; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2586 = 8'h12 == bh_iodex ? branch_target_buffer_18 : _GEN_2585; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2587 = 8'h13 == bh_iodex ? branch_target_buffer_19 : _GEN_2586; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2588 = 8'h14 == bh_iodex ? branch_target_buffer_20 : _GEN_2587; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2589 = 8'h15 == bh_iodex ? branch_target_buffer_21 : _GEN_2588; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2590 = 8'h16 == bh_iodex ? branch_target_buffer_22 : _GEN_2589; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2591 = 8'h17 == bh_iodex ? branch_target_buffer_23 : _GEN_2590; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2592 = 8'h18 == bh_iodex ? branch_target_buffer_24 : _GEN_2591; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2593 = 8'h19 == bh_iodex ? branch_target_buffer_25 : _GEN_2592; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2594 = 8'h1a == bh_iodex ? branch_target_buffer_26 : _GEN_2593; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2595 = 8'h1b == bh_iodex ? branch_target_buffer_27 : _GEN_2594; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2596 = 8'h1c == bh_iodex ? branch_target_buffer_28 : _GEN_2595; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2597 = 8'h1d == bh_iodex ? branch_target_buffer_29 : _GEN_2596; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2598 = 8'h1e == bh_iodex ? branch_target_buffer_30 : _GEN_2597; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2599 = 8'h1f == bh_iodex ? branch_target_buffer_31 : _GEN_2598; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2600 = 8'h20 == bh_iodex ? branch_target_buffer_32 : _GEN_2599; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2601 = 8'h21 == bh_iodex ? branch_target_buffer_33 : _GEN_2600; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2602 = 8'h22 == bh_iodex ? branch_target_buffer_34 : _GEN_2601; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2603 = 8'h23 == bh_iodex ? branch_target_buffer_35 : _GEN_2602; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2604 = 8'h24 == bh_iodex ? branch_target_buffer_36 : _GEN_2603; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2605 = 8'h25 == bh_iodex ? branch_target_buffer_37 : _GEN_2604; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2606 = 8'h26 == bh_iodex ? branch_target_buffer_38 : _GEN_2605; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2607 = 8'h27 == bh_iodex ? branch_target_buffer_39 : _GEN_2606; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2608 = 8'h28 == bh_iodex ? branch_target_buffer_40 : _GEN_2607; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2609 = 8'h29 == bh_iodex ? branch_target_buffer_41 : _GEN_2608; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2610 = 8'h2a == bh_iodex ? branch_target_buffer_42 : _GEN_2609; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2611 = 8'h2b == bh_iodex ? branch_target_buffer_43 : _GEN_2610; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2612 = 8'h2c == bh_iodex ? branch_target_buffer_44 : _GEN_2611; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2613 = 8'h2d == bh_iodex ? branch_target_buffer_45 : _GEN_2612; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2614 = 8'h2e == bh_iodex ? branch_target_buffer_46 : _GEN_2613; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2615 = 8'h2f == bh_iodex ? branch_target_buffer_47 : _GEN_2614; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2616 = 8'h30 == bh_iodex ? branch_target_buffer_48 : _GEN_2615; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2617 = 8'h31 == bh_iodex ? branch_target_buffer_49 : _GEN_2616; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2618 = 8'h32 == bh_iodex ? branch_target_buffer_50 : _GEN_2617; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2619 = 8'h33 == bh_iodex ? branch_target_buffer_51 : _GEN_2618; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2620 = 8'h34 == bh_iodex ? branch_target_buffer_52 : _GEN_2619; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2621 = 8'h35 == bh_iodex ? branch_target_buffer_53 : _GEN_2620; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2622 = 8'h36 == bh_iodex ? branch_target_buffer_54 : _GEN_2621; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2623 = 8'h37 == bh_iodex ? branch_target_buffer_55 : _GEN_2622; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2624 = 8'h38 == bh_iodex ? branch_target_buffer_56 : _GEN_2623; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2625 = 8'h39 == bh_iodex ? branch_target_buffer_57 : _GEN_2624; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2626 = 8'h3a == bh_iodex ? branch_target_buffer_58 : _GEN_2625; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2627 = 8'h3b == bh_iodex ? branch_target_buffer_59 : _GEN_2626; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2628 = 8'h3c == bh_iodex ? branch_target_buffer_60 : _GEN_2627; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2629 = 8'h3d == bh_iodex ? branch_target_buffer_61 : _GEN_2628; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2630 = 8'h3e == bh_iodex ? branch_target_buffer_62 : _GEN_2629; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2631 = 8'h3f == bh_iodex ? branch_target_buffer_63 : _GEN_2630; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2632 = 8'h40 == bh_iodex ? branch_target_buffer_64 : _GEN_2631; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2633 = 8'h41 == bh_iodex ? branch_target_buffer_65 : _GEN_2632; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2634 = 8'h42 == bh_iodex ? branch_target_buffer_66 : _GEN_2633; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2635 = 8'h43 == bh_iodex ? branch_target_buffer_67 : _GEN_2634; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2636 = 8'h44 == bh_iodex ? branch_target_buffer_68 : _GEN_2635; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2637 = 8'h45 == bh_iodex ? branch_target_buffer_69 : _GEN_2636; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2638 = 8'h46 == bh_iodex ? branch_target_buffer_70 : _GEN_2637; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2639 = 8'h47 == bh_iodex ? branch_target_buffer_71 : _GEN_2638; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2640 = 8'h48 == bh_iodex ? branch_target_buffer_72 : _GEN_2639; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2641 = 8'h49 == bh_iodex ? branch_target_buffer_73 : _GEN_2640; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2642 = 8'h4a == bh_iodex ? branch_target_buffer_74 : _GEN_2641; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2643 = 8'h4b == bh_iodex ? branch_target_buffer_75 : _GEN_2642; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2644 = 8'h4c == bh_iodex ? branch_target_buffer_76 : _GEN_2643; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2645 = 8'h4d == bh_iodex ? branch_target_buffer_77 : _GEN_2644; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2646 = 8'h4e == bh_iodex ? branch_target_buffer_78 : _GEN_2645; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2647 = 8'h4f == bh_iodex ? branch_target_buffer_79 : _GEN_2646; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2648 = 8'h50 == bh_iodex ? branch_target_buffer_80 : _GEN_2647; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2649 = 8'h51 == bh_iodex ? branch_target_buffer_81 : _GEN_2648; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2650 = 8'h52 == bh_iodex ? branch_target_buffer_82 : _GEN_2649; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2651 = 8'h53 == bh_iodex ? branch_target_buffer_83 : _GEN_2650; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2652 = 8'h54 == bh_iodex ? branch_target_buffer_84 : _GEN_2651; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2653 = 8'h55 == bh_iodex ? branch_target_buffer_85 : _GEN_2652; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2654 = 8'h56 == bh_iodex ? branch_target_buffer_86 : _GEN_2653; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2655 = 8'h57 == bh_iodex ? branch_target_buffer_87 : _GEN_2654; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2656 = 8'h58 == bh_iodex ? branch_target_buffer_88 : _GEN_2655; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2657 = 8'h59 == bh_iodex ? branch_target_buffer_89 : _GEN_2656; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2658 = 8'h5a == bh_iodex ? branch_target_buffer_90 : _GEN_2657; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2659 = 8'h5b == bh_iodex ? branch_target_buffer_91 : _GEN_2658; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2660 = 8'h5c == bh_iodex ? branch_target_buffer_92 : _GEN_2659; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2661 = 8'h5d == bh_iodex ? branch_target_buffer_93 : _GEN_2660; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2662 = 8'h5e == bh_iodex ? branch_target_buffer_94 : _GEN_2661; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2663 = 8'h5f == bh_iodex ? branch_target_buffer_95 : _GEN_2662; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2664 = 8'h60 == bh_iodex ? branch_target_buffer_96 : _GEN_2663; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2665 = 8'h61 == bh_iodex ? branch_target_buffer_97 : _GEN_2664; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2666 = 8'h62 == bh_iodex ? branch_target_buffer_98 : _GEN_2665; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2667 = 8'h63 == bh_iodex ? branch_target_buffer_99 : _GEN_2666; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2668 = 8'h64 == bh_iodex ? branch_target_buffer_100 : _GEN_2667; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2669 = 8'h65 == bh_iodex ? branch_target_buffer_101 : _GEN_2668; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2670 = 8'h66 == bh_iodex ? branch_target_buffer_102 : _GEN_2669; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2671 = 8'h67 == bh_iodex ? branch_target_buffer_103 : _GEN_2670; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2672 = 8'h68 == bh_iodex ? branch_target_buffer_104 : _GEN_2671; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2673 = 8'h69 == bh_iodex ? branch_target_buffer_105 : _GEN_2672; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2674 = 8'h6a == bh_iodex ? branch_target_buffer_106 : _GEN_2673; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2675 = 8'h6b == bh_iodex ? branch_target_buffer_107 : _GEN_2674; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2676 = 8'h6c == bh_iodex ? branch_target_buffer_108 : _GEN_2675; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2677 = 8'h6d == bh_iodex ? branch_target_buffer_109 : _GEN_2676; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2678 = 8'h6e == bh_iodex ? branch_target_buffer_110 : _GEN_2677; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2679 = 8'h6f == bh_iodex ? branch_target_buffer_111 : _GEN_2678; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2680 = 8'h70 == bh_iodex ? branch_target_buffer_112 : _GEN_2679; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2681 = 8'h71 == bh_iodex ? branch_target_buffer_113 : _GEN_2680; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2682 = 8'h72 == bh_iodex ? branch_target_buffer_114 : _GEN_2681; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2683 = 8'h73 == bh_iodex ? branch_target_buffer_115 : _GEN_2682; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2684 = 8'h74 == bh_iodex ? branch_target_buffer_116 : _GEN_2683; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2685 = 8'h75 == bh_iodex ? branch_target_buffer_117 : _GEN_2684; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2686 = 8'h76 == bh_iodex ? branch_target_buffer_118 : _GEN_2685; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2687 = 8'h77 == bh_iodex ? branch_target_buffer_119 : _GEN_2686; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2688 = 8'h78 == bh_iodex ? branch_target_buffer_120 : _GEN_2687; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2689 = 8'h79 == bh_iodex ? branch_target_buffer_121 : _GEN_2688; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2690 = 8'h7a == bh_iodex ? branch_target_buffer_122 : _GEN_2689; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2691 = 8'h7b == bh_iodex ? branch_target_buffer_123 : _GEN_2690; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2692 = 8'h7c == bh_iodex ? branch_target_buffer_124 : _GEN_2691; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2693 = 8'h7d == bh_iodex ? branch_target_buffer_125 : _GEN_2692; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2694 = 8'h7e == bh_iodex ? branch_target_buffer_126 : _GEN_2693; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2695 = 8'h7f == bh_iodex ? branch_target_buffer_127 : _GEN_2694; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2696 = 8'h80 == bh_iodex ? branch_target_buffer_128 : _GEN_2695; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2697 = 8'h81 == bh_iodex ? branch_target_buffer_129 : _GEN_2696; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2698 = 8'h82 == bh_iodex ? branch_target_buffer_130 : _GEN_2697; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2699 = 8'h83 == bh_iodex ? branch_target_buffer_131 : _GEN_2698; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2700 = 8'h84 == bh_iodex ? branch_target_buffer_132 : _GEN_2699; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2701 = 8'h85 == bh_iodex ? branch_target_buffer_133 : _GEN_2700; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2702 = 8'h86 == bh_iodex ? branch_target_buffer_134 : _GEN_2701; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2703 = 8'h87 == bh_iodex ? branch_target_buffer_135 : _GEN_2702; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2704 = 8'h88 == bh_iodex ? branch_target_buffer_136 : _GEN_2703; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2705 = 8'h89 == bh_iodex ? branch_target_buffer_137 : _GEN_2704; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2706 = 8'h8a == bh_iodex ? branch_target_buffer_138 : _GEN_2705; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2707 = 8'h8b == bh_iodex ? branch_target_buffer_139 : _GEN_2706; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2708 = 8'h8c == bh_iodex ? branch_target_buffer_140 : _GEN_2707; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2709 = 8'h8d == bh_iodex ? branch_target_buffer_141 : _GEN_2708; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2710 = 8'h8e == bh_iodex ? branch_target_buffer_142 : _GEN_2709; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2711 = 8'h8f == bh_iodex ? branch_target_buffer_143 : _GEN_2710; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2712 = 8'h90 == bh_iodex ? branch_target_buffer_144 : _GEN_2711; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2713 = 8'h91 == bh_iodex ? branch_target_buffer_145 : _GEN_2712; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2714 = 8'h92 == bh_iodex ? branch_target_buffer_146 : _GEN_2713; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2715 = 8'h93 == bh_iodex ? branch_target_buffer_147 : _GEN_2714; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2716 = 8'h94 == bh_iodex ? branch_target_buffer_148 : _GEN_2715; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2717 = 8'h95 == bh_iodex ? branch_target_buffer_149 : _GEN_2716; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2718 = 8'h96 == bh_iodex ? branch_target_buffer_150 : _GEN_2717; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2719 = 8'h97 == bh_iodex ? branch_target_buffer_151 : _GEN_2718; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2720 = 8'h98 == bh_iodex ? branch_target_buffer_152 : _GEN_2719; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2721 = 8'h99 == bh_iodex ? branch_target_buffer_153 : _GEN_2720; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2722 = 8'h9a == bh_iodex ? branch_target_buffer_154 : _GEN_2721; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2723 = 8'h9b == bh_iodex ? branch_target_buffer_155 : _GEN_2722; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2724 = 8'h9c == bh_iodex ? branch_target_buffer_156 : _GEN_2723; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2725 = 8'h9d == bh_iodex ? branch_target_buffer_157 : _GEN_2724; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2726 = 8'h9e == bh_iodex ? branch_target_buffer_158 : _GEN_2725; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2727 = 8'h9f == bh_iodex ? branch_target_buffer_159 : _GEN_2726; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2728 = 8'ha0 == bh_iodex ? branch_target_buffer_160 : _GEN_2727; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2729 = 8'ha1 == bh_iodex ? branch_target_buffer_161 : _GEN_2728; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2730 = 8'ha2 == bh_iodex ? branch_target_buffer_162 : _GEN_2729; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2731 = 8'ha3 == bh_iodex ? branch_target_buffer_163 : _GEN_2730; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2732 = 8'ha4 == bh_iodex ? branch_target_buffer_164 : _GEN_2731; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2733 = 8'ha5 == bh_iodex ? branch_target_buffer_165 : _GEN_2732; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2734 = 8'ha6 == bh_iodex ? branch_target_buffer_166 : _GEN_2733; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2735 = 8'ha7 == bh_iodex ? branch_target_buffer_167 : _GEN_2734; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2736 = 8'ha8 == bh_iodex ? branch_target_buffer_168 : _GEN_2735; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2737 = 8'ha9 == bh_iodex ? branch_target_buffer_169 : _GEN_2736; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2738 = 8'haa == bh_iodex ? branch_target_buffer_170 : _GEN_2737; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2739 = 8'hab == bh_iodex ? branch_target_buffer_171 : _GEN_2738; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2740 = 8'hac == bh_iodex ? branch_target_buffer_172 : _GEN_2739; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2741 = 8'had == bh_iodex ? branch_target_buffer_173 : _GEN_2740; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2742 = 8'hae == bh_iodex ? branch_target_buffer_174 : _GEN_2741; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2743 = 8'haf == bh_iodex ? branch_target_buffer_175 : _GEN_2742; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2744 = 8'hb0 == bh_iodex ? branch_target_buffer_176 : _GEN_2743; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2745 = 8'hb1 == bh_iodex ? branch_target_buffer_177 : _GEN_2744; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2746 = 8'hb2 == bh_iodex ? branch_target_buffer_178 : _GEN_2745; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2747 = 8'hb3 == bh_iodex ? branch_target_buffer_179 : _GEN_2746; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2748 = 8'hb4 == bh_iodex ? branch_target_buffer_180 : _GEN_2747; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2749 = 8'hb5 == bh_iodex ? branch_target_buffer_181 : _GEN_2748; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2750 = 8'hb6 == bh_iodex ? branch_target_buffer_182 : _GEN_2749; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2751 = 8'hb7 == bh_iodex ? branch_target_buffer_183 : _GEN_2750; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2752 = 8'hb8 == bh_iodex ? branch_target_buffer_184 : _GEN_2751; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2753 = 8'hb9 == bh_iodex ? branch_target_buffer_185 : _GEN_2752; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2754 = 8'hba == bh_iodex ? branch_target_buffer_186 : _GEN_2753; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2755 = 8'hbb == bh_iodex ? branch_target_buffer_187 : _GEN_2754; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2756 = 8'hbc == bh_iodex ? branch_target_buffer_188 : _GEN_2755; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2757 = 8'hbd == bh_iodex ? branch_target_buffer_189 : _GEN_2756; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2758 = 8'hbe == bh_iodex ? branch_target_buffer_190 : _GEN_2757; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2759 = 8'hbf == bh_iodex ? branch_target_buffer_191 : _GEN_2758; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2760 = 8'hc0 == bh_iodex ? branch_target_buffer_192 : _GEN_2759; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2761 = 8'hc1 == bh_iodex ? branch_target_buffer_193 : _GEN_2760; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2762 = 8'hc2 == bh_iodex ? branch_target_buffer_194 : _GEN_2761; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2763 = 8'hc3 == bh_iodex ? branch_target_buffer_195 : _GEN_2762; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2764 = 8'hc4 == bh_iodex ? branch_target_buffer_196 : _GEN_2763; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2765 = 8'hc5 == bh_iodex ? branch_target_buffer_197 : _GEN_2764; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2766 = 8'hc6 == bh_iodex ? branch_target_buffer_198 : _GEN_2765; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2767 = 8'hc7 == bh_iodex ? branch_target_buffer_199 : _GEN_2766; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2768 = 8'hc8 == bh_iodex ? branch_target_buffer_200 : _GEN_2767; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2769 = 8'hc9 == bh_iodex ? branch_target_buffer_201 : _GEN_2768; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2770 = 8'hca == bh_iodex ? branch_target_buffer_202 : _GEN_2769; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2771 = 8'hcb == bh_iodex ? branch_target_buffer_203 : _GEN_2770; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2772 = 8'hcc == bh_iodex ? branch_target_buffer_204 : _GEN_2771; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2773 = 8'hcd == bh_iodex ? branch_target_buffer_205 : _GEN_2772; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2774 = 8'hce == bh_iodex ? branch_target_buffer_206 : _GEN_2773; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2775 = 8'hcf == bh_iodex ? branch_target_buffer_207 : _GEN_2774; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2776 = 8'hd0 == bh_iodex ? branch_target_buffer_208 : _GEN_2775; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2777 = 8'hd1 == bh_iodex ? branch_target_buffer_209 : _GEN_2776; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2778 = 8'hd2 == bh_iodex ? branch_target_buffer_210 : _GEN_2777; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2779 = 8'hd3 == bh_iodex ? branch_target_buffer_211 : _GEN_2778; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2780 = 8'hd4 == bh_iodex ? branch_target_buffer_212 : _GEN_2779; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2781 = 8'hd5 == bh_iodex ? branch_target_buffer_213 : _GEN_2780; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2782 = 8'hd6 == bh_iodex ? branch_target_buffer_214 : _GEN_2781; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2783 = 8'hd7 == bh_iodex ? branch_target_buffer_215 : _GEN_2782; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2784 = 8'hd8 == bh_iodex ? branch_target_buffer_216 : _GEN_2783; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2785 = 8'hd9 == bh_iodex ? branch_target_buffer_217 : _GEN_2784; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2786 = 8'hda == bh_iodex ? branch_target_buffer_218 : _GEN_2785; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2787 = 8'hdb == bh_iodex ? branch_target_buffer_219 : _GEN_2786; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2788 = 8'hdc == bh_iodex ? branch_target_buffer_220 : _GEN_2787; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2789 = 8'hdd == bh_iodex ? branch_target_buffer_221 : _GEN_2788; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2790 = 8'hde == bh_iodex ? branch_target_buffer_222 : _GEN_2789; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2791 = 8'hdf == bh_iodex ? branch_target_buffer_223 : _GEN_2790; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2792 = 8'he0 == bh_iodex ? branch_target_buffer_224 : _GEN_2791; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2793 = 8'he1 == bh_iodex ? branch_target_buffer_225 : _GEN_2792; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2794 = 8'he2 == bh_iodex ? branch_target_buffer_226 : _GEN_2793; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2795 = 8'he3 == bh_iodex ? branch_target_buffer_227 : _GEN_2794; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2796 = 8'he4 == bh_iodex ? branch_target_buffer_228 : _GEN_2795; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2797 = 8'he5 == bh_iodex ? branch_target_buffer_229 : _GEN_2796; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2798 = 8'he6 == bh_iodex ? branch_target_buffer_230 : _GEN_2797; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2799 = 8'he7 == bh_iodex ? branch_target_buffer_231 : _GEN_2798; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2800 = 8'he8 == bh_iodex ? branch_target_buffer_232 : _GEN_2799; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2801 = 8'he9 == bh_iodex ? branch_target_buffer_233 : _GEN_2800; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2802 = 8'hea == bh_iodex ? branch_target_buffer_234 : _GEN_2801; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2803 = 8'heb == bh_iodex ? branch_target_buffer_235 : _GEN_2802; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2804 = 8'hec == bh_iodex ? branch_target_buffer_236 : _GEN_2803; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2805 = 8'hed == bh_iodex ? branch_target_buffer_237 : _GEN_2804; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2806 = 8'hee == bh_iodex ? branch_target_buffer_238 : _GEN_2805; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2807 = 8'hef == bh_iodex ? branch_target_buffer_239 : _GEN_2806; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2808 = 8'hf0 == bh_iodex ? branch_target_buffer_240 : _GEN_2807; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2809 = 8'hf1 == bh_iodex ? branch_target_buffer_241 : _GEN_2808; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2810 = 8'hf2 == bh_iodex ? branch_target_buffer_242 : _GEN_2809; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2811 = 8'hf3 == bh_iodex ? branch_target_buffer_243 : _GEN_2810; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2812 = 8'hf4 == bh_iodex ? branch_target_buffer_244 : _GEN_2811; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2813 = 8'hf5 == bh_iodex ? branch_target_buffer_245 : _GEN_2812; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2814 = 8'hf6 == bh_iodex ? branch_target_buffer_246 : _GEN_2813; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2815 = 8'hf7 == bh_iodex ? branch_target_buffer_247 : _GEN_2814; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2816 = 8'hf8 == bh_iodex ? branch_target_buffer_248 : _GEN_2815; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2817 = 8'hf9 == bh_iodex ? branch_target_buffer_249 : _GEN_2816; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2818 = 8'hfa == bh_iodex ? branch_target_buffer_250 : _GEN_2817; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2819 = 8'hfb == bh_iodex ? branch_target_buffer_251 : _GEN_2818; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2820 = 8'hfc == bh_iodex ? branch_target_buffer_252 : _GEN_2819; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2821 = 8'hfd == bh_iodex ? branch_target_buffer_253 : _GEN_2820; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2822 = 8'hfe == bh_iodex ? branch_target_buffer_254 : _GEN_2821; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _GEN_2823 = 8'hff == bh_iodex ? branch_target_buffer_255 : _GEN_2822; // @[BP.scala 128:51 BP.scala 128:51]
  wire [31:0] _pred_target_T_3 = io_in_pc_io_reg_pc + 32'h4; // @[BP.scala 128:77]
  assign io_out_pred_flag = pt_flag ? _T_5 : _T_10; // @[BP.scala 114:19]
  assign io_out_pred_target = pred_flag & _GEN_2823 != 32'h0 ? _GEN_2823 : _pred_target_T_3; // @[BP.scala 128:27]
  always @(posedge clock) begin
    if (reset) begin // @[BP.scala 53:42]
      branch_history_0 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_0 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_0 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_1 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_1 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_1 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_2 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_2 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_2 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_3 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_3 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_3 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_4 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_4 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_4 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_5 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_5 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_5 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_6 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_6 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_6 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_7 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_7 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_7 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_8 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_8 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_8 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_9 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_9 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_9 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_10 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_10 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_10 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_11 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_11 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_11 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_12 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_12 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_12 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_13 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_13 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_13 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_14 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_14 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_14 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_15 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_15 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_15 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_16 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h10 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_16 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_16 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_17 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h11 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_17 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_17 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_18 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h12 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_18 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_18 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_19 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h13 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_19 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_19 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_20 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h14 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_20 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_20 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_21 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h15 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_21 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_21 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_22 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h16 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_22 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_22 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_23 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h17 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_23 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_23 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_24 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h18 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_24 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_24 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_25 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h19 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_25 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_25 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_26 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_26 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_26 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_27 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_27 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_27 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_28 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_28 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_28 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_29 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_29 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_29 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_30 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_30 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_30 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_31 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_31 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_31 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_32 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h20 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_32 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_32 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_33 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h21 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_33 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_33 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_34 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h22 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_34 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_34 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_35 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h23 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_35 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_35 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_36 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h24 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_36 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_36 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_37 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h25 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_37 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_37 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_38 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h26 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_38 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_38 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_39 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h27 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_39 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_39 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_40 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h28 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_40 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_40 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_41 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h29 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_41 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_41 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_42 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_42 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_42 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_43 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_43 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_43 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_44 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_44 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_44 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_45 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_45 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_45 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_46 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_46 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_46 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_47 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_47 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_47 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_48 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h30 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_48 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_48 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_49 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h31 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_49 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_49 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_50 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h32 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_50 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_50 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_51 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h33 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_51 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_51 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_52 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h34 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_52 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_52 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_53 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h35 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_53 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_53 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_54 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h36 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_54 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_54 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_55 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h37 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_55 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_55 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_56 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h38 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_56 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_56 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_57 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h39 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_57 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_57 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_58 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_58 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_58 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_59 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_59 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_59 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_60 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_60 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_60 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_61 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_61 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_61 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_62 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_62 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_62 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_63 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_63 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_63 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_64 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h40 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_64 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_64 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_65 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h41 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_65 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_65 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_66 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h42 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_66 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_66 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_67 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h43 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_67 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_67 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_68 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h44 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_68 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_68 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_69 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h45 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_69 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_69 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_70 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h46 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_70 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_70 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_71 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h47 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_71 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_71 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_72 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h48 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_72 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_72 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_73 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h49 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_73 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_73 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_74 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_74 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_74 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_75 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_75 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_75 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_76 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_76 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_76 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_77 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_77 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_77 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_78 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_78 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_78 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_79 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_79 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_79 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_80 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h50 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_80 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_80 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_81 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h51 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_81 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_81 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_82 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h52 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_82 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_82 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_83 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h53 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_83 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_83 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_84 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h54 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_84 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_84 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_85 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h55 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_85 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_85 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_86 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h56 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_86 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_86 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_87 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h57 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_87 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_87 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_88 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h58 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_88 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_88 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_89 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h59 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_89 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_89 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_90 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_90 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_90 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_91 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_91 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_91 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_92 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_92 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_92 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_93 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_93 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_93 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_94 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_94 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_94 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_95 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_95 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_95 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_96 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h60 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_96 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_96 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_97 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h61 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_97 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_97 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_98 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h62 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_98 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_98 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_99 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h63 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_99 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_99 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_100 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h64 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_100 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_100 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_101 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h65 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_101 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_101 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_102 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h66 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_102 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_102 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_103 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h67 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_103 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_103 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_104 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h68 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_104 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_104 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_105 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h69 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_105 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_105 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_106 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_106 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_106 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_107 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_107 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_107 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_108 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_108 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_108 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_109 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_109 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_109 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_110 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_110 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_110 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_111 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_111 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_111 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_112 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h70 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_112 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_112 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_113 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h71 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_113 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_113 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_114 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h72 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_114 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_114 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_115 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h73 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_115 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_115 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_116 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h74 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_116 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_116 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_117 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h75 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_117 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_117 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_118 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h76 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_118 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_118 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_119 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h77 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_119 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_119 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_120 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h78 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_120 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_120 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_121 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h79 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_121 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_121 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_122 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_122 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_122 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_123 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_123 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_123 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_124 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_124 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_124 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_125 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_125 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_125 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_126 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_126 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_126 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_127 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_127 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_127 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_128 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h80 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_128 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_128 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_129 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h81 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_129 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_129 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_130 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h82 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_130 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_130 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_131 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h83 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_131 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_131 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_132 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h84 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_132 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_132 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_133 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h85 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_133 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_133 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_134 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h86 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_134 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_134 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_135 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h87 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_135 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_135 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_136 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h88 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_136 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_136 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_137 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h89 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_137 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_137 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_138 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_138 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_138 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_139 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_139 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_139 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_140 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_140 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_140 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_141 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_141 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_141 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_142 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_142 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_142 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_143 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_143 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_143 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_144 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h90 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_144 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_144 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_145 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h91 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_145 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_145 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_146 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h92 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_146 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_146 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_147 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h93 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_147 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_147 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_148 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h94 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_148 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_148 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_149 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h95 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_149 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_149 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_150 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h96 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_150 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_150 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_151 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h97 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_151 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_151 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_152 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h98 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_152 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_152 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_153 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h99 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_153 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_153 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_154 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9a == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_154 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_154 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_155 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9b == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_155 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_155 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_156 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9c == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_156 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_156 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_157 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9d == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_157 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_157 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_158 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9e == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_158 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_158 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_159 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9f == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_159 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_159 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_160 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_160 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_160 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_161 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_161 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_161 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_162 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_162 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_162 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_163 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_163 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_163 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_164 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_164 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_164 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_165 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_165 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_165 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_166 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_166 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_166 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_167 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_167 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_167 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_168 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_168 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_168 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_169 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_169 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_169 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_170 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'haa == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_170 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_170 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_171 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hab == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_171 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_171 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_172 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hac == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_172 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_172 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_173 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'had == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_173 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_173 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_174 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hae == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_174 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_174 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_175 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'haf == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_175 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_175 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_176 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_176 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_176 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_177 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_177 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_177 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_178 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_178 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_178 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_179 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_179 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_179 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_180 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_180 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_180 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_181 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_181 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_181 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_182 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_182 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_182 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_183 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_183 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_183 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_184 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_184 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_184 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_185 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_185 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_185 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_186 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hba == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_186 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_186 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_187 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_187 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_187 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_188 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbc == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_188 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_188 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_189 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbd == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_189 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_189 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_190 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbe == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_190 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_190 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_191 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbf == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_191 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_191 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_192 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_192 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_192 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_193 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_193 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_193 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_194 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_194 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_194 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_195 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_195 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_195 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_196 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_196 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_196 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_197 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_197 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_197 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_198 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_198 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_198 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_199 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_199 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_199 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_200 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_200 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_200 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_201 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_201 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_201 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_202 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hca == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_202 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_202 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_203 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_203 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_203 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_204 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcc == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_204 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_204 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_205 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcd == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_205 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_205 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_206 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hce == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_206 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_206 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_207 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcf == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_207 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_207 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_208 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_208 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_208 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_209 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_209 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_209 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_210 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_210 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_210 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_211 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_211 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_211 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_212 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_212 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_212 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_213 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_213 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_213 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_214 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_214 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_214 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_215 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_215 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_215 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_216 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_216 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_216 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_217 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_217 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_217 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_218 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hda == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_218 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_218 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_219 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_219 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_219 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_220 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdc == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_220 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_220 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_221 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdd == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_221 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_221 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_222 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hde == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_222 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_222 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_223 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdf == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_223 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_223 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_224 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_224 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_224 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_225 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_225 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_225 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_226 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_226 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_226 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_227 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_227 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_227 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_228 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_228 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_228 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_229 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_229 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_229 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_230 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_230 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_230 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_231 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_231 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_231 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_232 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_232 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_232 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_233 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_233 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_233 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_234 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hea == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_234 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_234 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_235 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'heb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_235 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_235 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_236 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hec == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_236 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_236 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_237 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hed == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_237 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_237 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_238 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hee == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_238 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_238 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_239 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hef == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_239 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_239 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_240 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf0 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_240 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_240 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_241 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf1 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_241 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_241 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_242 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf2 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_242 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_242 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_243 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf3 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_243 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_243 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_244 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf4 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_244 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_244 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_245 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf5 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_245 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_245 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_246 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf6 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_246 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_246 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_247 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf7 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_247 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_247 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_248 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf8 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_248 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_248 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_249 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf9 == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_249 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_249 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_250 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfa == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_250 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_250 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_251 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfb == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_251 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_251 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_252 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfc == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_252 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_252 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_253 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfd == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_253 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_253 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_254 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfe == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_254 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_254 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 53:42]
      branch_history_255 <= 8'h0; // @[BP.scala 53:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hff == ex_bh_iodex) begin // @[BP.scala 91:37]
        if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
          branch_history_255 <= _new_bh_value_T_2; // @[BP.scala 90:22]
        end else begin
          branch_history_255 <= shifted_bh; // @[BP.scala 87:21]
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_0 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_0 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_0 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_1 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_1 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_1 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_2 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_2 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_2 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_3 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_3 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_3 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_4 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_4 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_4 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_5 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_5 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_5 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_6 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_6 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_6 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_7 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_7 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_7 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_8 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_8 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_8 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_9 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_9 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_9 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_10 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_10 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_10 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_11 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_11 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_11 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_12 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_12 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_12 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_13 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_13 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_13 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_14 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_14 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_14 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_15 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_15 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_15 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_16 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h10 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_16 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_16 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_17 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h11 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_17 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_17 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_18 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h12 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_18 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_18 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_19 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h13 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_19 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_19 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_20 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h14 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_20 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_20 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_21 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h15 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_21 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_21 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_22 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h16 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_22 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_22 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_23 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h17 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_23 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_23 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_24 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h18 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_24 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_24 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_25 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h19 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_25 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_25 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_26 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_26 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_26 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_27 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_27 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_27 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_28 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_28 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_28 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_29 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_29 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_29 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_30 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_30 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_30 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_31 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h1f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_31 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_31 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_32 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h20 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_32 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_32 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_33 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h21 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_33 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_33 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_34 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h22 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_34 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_34 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_35 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h23 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_35 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_35 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_36 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h24 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_36 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_36 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_37 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h25 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_37 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_37 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_38 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h26 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_38 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_38 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_39 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h27 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_39 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_39 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_40 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h28 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_40 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_40 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_41 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h29 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_41 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_41 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_42 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_42 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_42 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_43 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_43 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_43 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_44 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_44 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_44 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_45 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_45 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_45 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_46 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_46 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_46 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_47 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h2f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_47 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_47 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_48 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h30 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_48 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_48 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_49 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h31 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_49 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_49 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_50 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h32 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_50 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_50 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_51 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h33 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_51 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_51 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_52 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h34 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_52 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_52 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_53 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h35 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_53 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_53 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_54 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h36 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_54 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_54 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_55 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h37 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_55 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_55 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_56 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h38 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_56 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_56 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_57 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h39 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_57 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_57 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_58 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_58 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_58 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_59 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_59 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_59 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_60 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_60 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_60 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_61 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_61 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_61 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_62 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_62 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_62 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_63 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h3f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_63 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_63 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_64 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h40 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_64 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_64 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_65 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h41 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_65 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_65 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_66 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h42 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_66 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_66 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_67 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h43 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_67 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_67 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_68 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h44 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_68 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_68 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_69 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h45 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_69 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_69 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_70 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h46 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_70 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_70 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_71 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h47 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_71 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_71 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_72 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h48 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_72 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_72 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_73 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h49 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_73 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_73 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_74 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_74 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_74 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_75 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_75 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_75 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_76 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_76 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_76 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_77 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_77 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_77 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_78 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_78 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_78 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_79 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h4f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_79 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_79 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_80 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h50 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_80 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_80 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_81 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h51 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_81 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_81 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_82 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h52 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_82 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_82 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_83 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h53 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_83 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_83 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_84 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h54 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_84 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_84 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_85 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h55 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_85 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_85 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_86 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h56 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_86 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_86 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_87 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h57 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_87 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_87 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_88 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h58 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_88 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_88 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_89 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h59 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_89 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_89 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_90 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_90 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_90 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_91 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_91 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_91 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_92 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_92 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_92 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_93 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_93 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_93 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_94 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_94 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_94 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_95 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h5f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_95 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_95 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_96 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h60 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_96 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_96 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_97 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h61 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_97 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_97 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_98 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h62 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_98 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_98 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_99 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h63 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_99 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_99 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_100 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h64 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_100 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_100 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_101 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h65 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_101 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_101 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_102 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h66 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_102 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_102 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_103 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h67 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_103 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_103 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_104 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h68 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_104 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_104 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_105 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h69 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_105 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_105 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_106 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_106 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_106 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_107 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_107 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_107 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_108 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_108 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_108 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_109 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_109 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_109 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_110 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_110 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_110 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_111 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h6f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_111 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_111 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_112 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h70 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_112 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_112 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_113 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h71 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_113 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_113 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_114 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h72 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_114 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_114 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_115 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h73 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_115 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_115 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_116 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h74 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_116 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_116 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_117 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h75 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_117 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_117 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_118 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h76 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_118 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_118 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_119 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h77 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_119 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_119 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_120 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h78 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_120 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_120 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_121 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h79 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_121 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_121 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_122 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_122 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_122 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_123 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_123 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_123 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_124 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_124 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_124 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_125 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_125 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_125 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_126 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_126 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_126 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_127 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h7f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_127 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_127 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_128 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h80 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_128 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_128 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_129 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h81 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_129 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_129 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_130 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h82 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_130 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_130 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_131 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h83 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_131 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_131 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_132 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h84 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_132 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_132 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_133 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h85 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_133 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_133 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_134 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h86 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_134 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_134 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_135 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h87 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_135 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_135 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_136 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h88 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_136 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_136 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_137 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h89 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_137 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_137 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_138 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_138 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_138 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_139 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_139 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_139 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_140 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_140 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_140 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_141 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_141 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_141 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_142 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_142 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_142 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_143 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h8f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_143 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_143 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_144 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h90 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_144 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_144 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_145 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h91 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_145 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_145 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_146 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h92 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_146 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_146 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_147 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h93 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_147 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_147 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_148 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h94 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_148 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_148 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_149 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h95 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_149 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_149 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_150 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h96 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_150 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_150 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_151 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h97 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_151 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_151 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_152 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h98 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_152 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_152 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_153 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h99 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_153 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_153 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_154 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9a == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_154 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_154 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_155 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9b == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_155 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_155 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_156 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9c == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_156 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_156 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_157 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9d == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_157 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_157 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_158 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9e == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_158 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_158 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_159 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'h9f == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_159 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_159 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_160 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_160 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_160 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_161 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_161 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_161 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_162 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_162 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_162 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_163 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_163 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_163 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_164 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_164 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_164 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_165 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_165 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_165 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_166 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_166 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_166 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_167 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_167 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_167 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_168 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_168 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_168 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_169 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'ha9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_169 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_169 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_170 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'haa == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_170 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_170 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_171 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hab == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_171 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_171 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_172 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hac == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_172 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_172 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_173 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'had == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_173 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_173 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_174 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hae == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_174 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_174 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_175 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'haf == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_175 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_175 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_176 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_176 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_176 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_177 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_177 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_177 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_178 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_178 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_178 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_179 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_179 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_179 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_180 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_180 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_180 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_181 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_181 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_181 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_182 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_182 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_182 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_183 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_183 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_183 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_184 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_184 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_184 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_185 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hb9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_185 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_185 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_186 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hba == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_186 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_186 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_187 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_187 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_187 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_188 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbc == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_188 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_188 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_189 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbd == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_189 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_189 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_190 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbe == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_190 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_190 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_191 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hbf == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_191 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_191 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_192 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_192 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_192 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_193 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_193 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_193 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_194 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_194 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_194 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_195 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_195 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_195 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_196 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_196 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_196 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_197 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_197 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_197 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_198 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_198 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_198 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_199 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_199 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_199 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_200 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_200 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_200 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_201 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hc9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_201 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_201 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_202 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hca == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_202 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_202 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_203 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_203 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_203 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_204 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcc == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_204 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_204 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_205 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcd == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_205 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_205 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_206 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hce == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_206 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_206 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_207 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hcf == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_207 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_207 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_208 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_208 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_208 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_209 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_209 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_209 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_210 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_210 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_210 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_211 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_211 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_211 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_212 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_212 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_212 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_213 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_213 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_213 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_214 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_214 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_214 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_215 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_215 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_215 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_216 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_216 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_216 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_217 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hd9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_217 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_217 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_218 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hda == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_218 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_218 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_219 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_219 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_219 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_220 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdc == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_220 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_220 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_221 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdd == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_221 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_221 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_222 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hde == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_222 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_222 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_223 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hdf == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_223 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_223 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_224 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_224 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_224 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_225 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_225 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_225 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_226 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_226 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_226 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_227 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_227 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_227 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_228 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_228 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_228 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_229 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_229 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_229 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_230 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_230 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_230 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_231 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_231 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_231 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_232 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_232 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_232 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_233 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'he9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_233 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_233 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_234 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hea == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_234 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_234 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_235 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'heb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_235 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_235 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_236 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hec == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_236 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_236 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_237 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hed == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_237 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_237 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_238 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hee == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_238 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_238 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_239 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hef == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_239 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_239 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_240 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf0 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_240 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_240 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_241 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf1 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_241 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_241 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_242 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf2 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_242 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_242 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_243 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf3 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_243 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_243 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_244 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf4 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_244 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_244 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_245 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf5 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_245 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_245 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_246 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf6 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_246 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_246 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_247 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf7 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_247 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_247 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_248 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf8 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_248 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_248 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_249 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hf9 == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_249 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_249 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_250 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfa == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_250 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_250 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_251 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfb == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_251 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_251 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_252 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfc == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_252 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_252 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_253 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfd == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_253 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_253 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_254 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hfe == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_254 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_254 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 54:42]
      pattern_table_255 <= 2'h1; // @[BP.scala 54:42]
    end else if (io_in_ex_io_br_io_pt_flag) begin // @[BP.scala 88:21]
      if (8'hff == new_bh_value) begin // @[BP.scala 92:37]
        if (_pattern_table_T) begin // @[Conditional.scala 40:58]
          pattern_table_255 <= _pattern_table_new_state_T; // @[BP.scala 79:33]
        end else begin
          pattern_table_255 <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_0 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_0 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_0 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_1 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_1 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_1 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_2 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_2 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_2 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_3 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_3 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_3 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_4 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_4 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_4 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_5 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_5 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_5 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_6 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_6 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_6 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_7 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_7 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_7 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_8 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_8 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_8 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_9 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_9 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_9 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_10 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_10 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_10 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_11 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_11 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_11 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_12 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_12 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_12 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_13 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_13 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_13 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_14 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_14 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_14 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_15 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_15 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_15 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_16 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h10 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_16 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_16 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_17 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h11 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_17 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_17 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_18 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h12 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_18 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_18 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_19 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h13 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_19 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_19 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_20 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h14 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_20 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_20 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_21 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h15 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_21 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_21 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_22 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h16 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_22 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_22 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_23 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h17 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_23 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_23 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_24 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h18 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_24 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_24 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_25 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h19 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_25 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_25 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_26 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_26 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_26 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_27 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_27 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_27 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_28 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_28 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_28 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_29 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_29 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_29 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_30 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_30 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_30 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_31 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h1f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_31 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_31 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_32 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h20 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_32 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_32 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_33 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h21 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_33 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_33 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_34 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h22 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_34 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_34 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_35 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h23 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_35 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_35 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_36 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h24 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_36 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_36 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_37 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h25 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_37 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_37 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_38 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h26 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_38 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_38 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_39 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h27 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_39 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_39 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_40 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h28 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_40 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_40 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_41 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h29 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_41 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_41 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_42 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_42 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_42 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_43 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_43 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_43 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_44 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_44 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_44 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_45 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_45 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_45 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_46 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_46 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_46 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_47 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h2f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_47 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_47 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_48 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h30 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_48 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_48 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_49 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h31 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_49 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_49 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_50 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h32 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_50 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_50 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_51 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h33 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_51 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_51 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_52 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h34 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_52 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_52 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_53 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h35 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_53 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_53 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_54 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h36 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_54 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_54 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_55 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h37 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_55 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_55 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_56 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h38 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_56 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_56 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_57 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h39 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_57 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_57 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_58 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_58 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_58 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_59 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_59 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_59 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_60 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_60 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_60 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_61 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_61 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_61 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_62 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_62 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_62 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_63 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h3f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_63 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_63 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_64 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h40 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_64 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_64 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_65 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h41 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_65 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_65 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_66 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h42 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_66 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_66 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_67 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h43 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_67 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_67 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_68 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h44 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_68 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_68 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_69 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h45 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_69 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_69 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_70 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h46 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_70 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_70 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_71 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h47 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_71 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_71 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_72 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h48 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_72 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_72 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_73 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h49 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_73 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_73 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_74 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_74 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_74 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_75 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_75 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_75 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_76 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_76 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_76 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_77 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_77 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_77 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_78 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_78 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_78 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_79 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h4f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_79 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_79 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_80 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h50 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_80 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_80 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_81 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h51 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_81 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_81 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_82 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h52 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_82 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_82 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_83 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h53 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_83 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_83 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_84 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h54 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_84 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_84 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_85 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h55 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_85 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_85 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_86 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h56 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_86 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_86 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_87 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h57 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_87 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_87 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_88 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h58 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_88 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_88 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_89 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h59 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_89 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_89 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_90 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_90 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_90 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_91 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_91 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_91 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_92 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_92 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_92 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_93 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_93 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_93 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_94 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_94 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_94 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_95 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h5f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_95 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_95 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_96 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h60 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_96 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_96 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_97 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h61 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_97 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_97 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_98 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h62 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_98 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_98 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_99 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h63 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_99 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_99 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_100 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h64 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_100 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_100 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_101 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h65 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_101 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_101 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_102 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h66 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_102 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_102 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_103 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h67 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_103 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_103 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_104 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h68 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_104 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_104 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_105 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h69 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_105 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_105 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_106 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_106 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_106 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_107 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_107 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_107 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_108 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_108 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_108 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_109 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_109 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_109 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_110 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_110 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_110 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_111 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h6f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_111 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_111 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_112 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h70 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_112 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_112 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_113 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h71 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_113 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_113 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_114 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h72 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_114 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_114 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_115 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h73 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_115 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_115 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_116 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h74 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_116 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_116 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_117 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h75 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_117 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_117 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_118 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h76 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_118 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_118 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_119 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h77 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_119 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_119 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_120 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h78 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_120 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_120 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_121 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h79 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_121 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_121 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_122 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_122 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_122 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_123 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_123 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_123 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_124 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_124 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_124 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_125 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_125 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_125 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_126 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_126 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_126 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_127 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h7f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_127 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_127 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_128 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h80 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_128 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_128 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_129 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h81 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_129 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_129 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_130 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h82 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_130 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_130 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_131 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h83 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_131 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_131 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_132 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h84 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_132 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_132 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_133 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h85 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_133 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_133 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_134 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h86 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_134 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_134 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_135 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h87 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_135 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_135 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_136 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h88 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_136 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_136 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_137 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h89 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_137 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_137 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_138 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_138 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_138 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_139 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_139 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_139 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_140 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_140 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_140 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_141 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_141 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_141 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_142 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_142 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_142 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_143 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h8f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_143 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_143 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_144 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h90 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_144 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_144 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_145 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h91 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_145 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_145 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_146 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h92 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_146 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_146 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_147 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h93 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_147 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_147 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_148 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h94 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_148 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_148 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_149 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h95 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_149 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_149 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_150 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h96 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_150 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_150 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_151 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h97 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_151 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_151 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_152 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h98 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_152 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_152 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_153 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h99 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_153 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_153 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_154 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9a == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_154 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_154 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_155 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9b == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_155 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_155 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_156 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9c == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_156 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_156 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_157 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9d == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_157 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_157 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_158 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9e == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_158 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_158 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_159 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'h9f == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_159 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_159 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_160 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_160 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_160 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_161 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_161 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_161 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_162 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_162 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_162 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_163 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_163 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_163 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_164 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_164 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_164 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_165 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_165 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_165 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_166 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_166 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_166 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_167 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_167 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_167 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_168 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_168 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_168 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_169 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'ha9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_169 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_169 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_170 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'haa == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_170 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_170 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_171 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hab == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_171 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_171 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_172 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hac == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_172 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_172 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_173 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'had == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_173 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_173 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_174 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hae == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_174 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_174 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_175 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'haf == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_175 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_175 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_176 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_176 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_176 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_177 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_177 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_177 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_178 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_178 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_178 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_179 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_179 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_179 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_180 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_180 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_180 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_181 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_181 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_181 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_182 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_182 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_182 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_183 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_183 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_183 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_184 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_184 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_184 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_185 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hb9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_185 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_185 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_186 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hba == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_186 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_186 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_187 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hbb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_187 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_187 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_188 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hbc == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_188 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_188 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_189 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hbd == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_189 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_189 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_190 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hbe == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_190 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_190 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_191 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hbf == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_191 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_191 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_192 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_192 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_192 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_193 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_193 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_193 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_194 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_194 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_194 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_195 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_195 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_195 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_196 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_196 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_196 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_197 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_197 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_197 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_198 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_198 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_198 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_199 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_199 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_199 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_200 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_200 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_200 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_201 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hc9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_201 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_201 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_202 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hca == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_202 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_202 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_203 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hcb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_203 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_203 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_204 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hcc == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_204 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_204 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_205 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hcd == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_205 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_205 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_206 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hce == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_206 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_206 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_207 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hcf == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_207 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_207 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_208 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_208 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_208 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_209 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_209 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_209 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_210 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_210 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_210 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_211 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_211 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_211 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_212 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_212 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_212 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_213 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_213 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_213 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_214 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_214 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_214 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_215 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_215 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_215 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_216 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_216 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_216 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_217 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hd9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_217 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_217 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_218 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hda == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_218 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_218 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_219 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hdb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_219 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_219 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_220 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hdc == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_220 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_220 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_221 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hdd == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_221 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_221 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_222 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hde == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_222 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_222 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_223 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hdf == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_223 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_223 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_224 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_224 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_224 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_225 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_225 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_225 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_226 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_226 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_226 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_227 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_227 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_227 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_228 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_228 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_228 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_229 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_229 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_229 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_230 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_230 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_230 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_231 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_231 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_231 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_232 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_232 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_232 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_233 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'he9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_233 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_233 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_234 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hea == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_234 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_234 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_235 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'heb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_235 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_235 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_236 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hec == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_236 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_236 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_237 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hed == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_237 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_237 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_238 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hee == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_238 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_238 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_239 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hef == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_239 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_239 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_240 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf0 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_240 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_240 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_241 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf1 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_241 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_241 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_242 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf2 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_242 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_242 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_243 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf3 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_243 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_243 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_244 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf4 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_244 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_244 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_245 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf5 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_245 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_245 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_246 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf6 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_246 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_246 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_247 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf7 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_247 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_247 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_248 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf8 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_248 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_248 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_249 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hf9 == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_249 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_249 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_250 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hfa == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_250 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_250 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_251 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hfb == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_251 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_251 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_252 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hfc == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_252 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_252 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_253 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hfd == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_253 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_253 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_254 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hfe == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_254 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_254 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
    if (reset) begin // @[BP.scala 55:42]
      branch_target_buffer_255 <= 32'h0; // @[BP.scala 55:42]
    end else if (io_in_ex_io_br_io_br_flag | io_in_ex_io_alu_io_jump_flag) begin // @[BP.scala 94:32]
      if (8'hff == ex_bh_iodex) begin // @[BP.scala 96:43]
        if (io_in_ex_io_br_io_br_flag) begin // @[BP.scala 96:49]
          branch_target_buffer_255 <= io_in_ex_io_br_io_br_target;
        end else begin
          branch_target_buffer_255 <= io_in_ex_io_alu_io_alu_out;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  branch_history_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  branch_history_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  branch_history_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  branch_history_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  branch_history_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  branch_history_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  branch_history_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  branch_history_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  branch_history_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  branch_history_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  branch_history_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  branch_history_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  branch_history_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  branch_history_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  branch_history_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  branch_history_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  branch_history_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  branch_history_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  branch_history_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  branch_history_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  branch_history_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  branch_history_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  branch_history_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  branch_history_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  branch_history_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  branch_history_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  branch_history_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  branch_history_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  branch_history_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  branch_history_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  branch_history_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  branch_history_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  branch_history_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  branch_history_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  branch_history_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  branch_history_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  branch_history_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  branch_history_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  branch_history_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  branch_history_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  branch_history_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  branch_history_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  branch_history_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  branch_history_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  branch_history_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  branch_history_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  branch_history_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  branch_history_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  branch_history_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  branch_history_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  branch_history_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  branch_history_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  branch_history_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  branch_history_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  branch_history_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  branch_history_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  branch_history_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  branch_history_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  branch_history_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  branch_history_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  branch_history_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  branch_history_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  branch_history_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  branch_history_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  branch_history_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  branch_history_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  branch_history_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  branch_history_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  branch_history_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  branch_history_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  branch_history_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  branch_history_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  branch_history_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  branch_history_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  branch_history_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  branch_history_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  branch_history_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  branch_history_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  branch_history_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  branch_history_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  branch_history_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  branch_history_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  branch_history_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  branch_history_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  branch_history_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  branch_history_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  branch_history_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  branch_history_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  branch_history_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  branch_history_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  branch_history_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  branch_history_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  branch_history_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  branch_history_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  branch_history_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  branch_history_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  branch_history_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  branch_history_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  branch_history_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  branch_history_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  branch_history_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  branch_history_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  branch_history_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  branch_history_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  branch_history_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  branch_history_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  branch_history_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  branch_history_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  branch_history_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  branch_history_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  branch_history_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  branch_history_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  branch_history_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  branch_history_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  branch_history_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  branch_history_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  branch_history_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  branch_history_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  branch_history_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  branch_history_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  branch_history_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  branch_history_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  branch_history_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  branch_history_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  branch_history_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  branch_history_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  branch_history_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  branch_history_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  branch_history_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  branch_history_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  branch_history_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  branch_history_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  branch_history_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  branch_history_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  branch_history_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  branch_history_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  branch_history_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  branch_history_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  branch_history_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  branch_history_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  branch_history_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  branch_history_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  branch_history_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  branch_history_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  branch_history_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  branch_history_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  branch_history_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  branch_history_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  branch_history_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  branch_history_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  branch_history_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  branch_history_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  branch_history_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  branch_history_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  branch_history_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  branch_history_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  branch_history_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  branch_history_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  branch_history_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  branch_history_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  branch_history_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  branch_history_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  branch_history_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  branch_history_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  branch_history_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  branch_history_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  branch_history_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  branch_history_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  branch_history_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  branch_history_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  branch_history_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  branch_history_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  branch_history_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  branch_history_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  branch_history_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  branch_history_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  branch_history_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  branch_history_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  branch_history_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  branch_history_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  branch_history_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  branch_history_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  branch_history_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  branch_history_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  branch_history_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  branch_history_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  branch_history_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  branch_history_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  branch_history_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  branch_history_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  branch_history_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  branch_history_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  branch_history_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  branch_history_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  branch_history_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  branch_history_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  branch_history_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  branch_history_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  branch_history_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  branch_history_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  branch_history_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  branch_history_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  branch_history_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  branch_history_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  branch_history_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  branch_history_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  branch_history_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  branch_history_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  branch_history_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  branch_history_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  branch_history_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  branch_history_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  branch_history_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  branch_history_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  branch_history_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  branch_history_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  branch_history_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  branch_history_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  branch_history_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  branch_history_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  branch_history_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  branch_history_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  branch_history_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  branch_history_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  branch_history_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  branch_history_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  branch_history_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  branch_history_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  branch_history_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  branch_history_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  branch_history_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  branch_history_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  branch_history_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  branch_history_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  branch_history_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  branch_history_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  branch_history_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  branch_history_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  branch_history_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  branch_history_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  branch_history_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  branch_history_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  branch_history_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  branch_history_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  branch_history_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  branch_history_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  branch_history_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  branch_history_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  branch_history_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  branch_history_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  branch_history_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  branch_history_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  branch_history_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  branch_history_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  branch_history_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  branch_history_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  pattern_table_0 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pattern_table_1 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pattern_table_2 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pattern_table_3 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pattern_table_4 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pattern_table_5 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pattern_table_6 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pattern_table_7 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pattern_table_8 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pattern_table_9 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pattern_table_10 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pattern_table_11 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pattern_table_12 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pattern_table_13 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pattern_table_14 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pattern_table_15 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pattern_table_16 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pattern_table_17 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pattern_table_18 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pattern_table_19 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pattern_table_20 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pattern_table_21 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pattern_table_22 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pattern_table_23 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pattern_table_24 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pattern_table_25 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pattern_table_26 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pattern_table_27 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pattern_table_28 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pattern_table_29 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pattern_table_30 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pattern_table_31 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pattern_table_32 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pattern_table_33 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pattern_table_34 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pattern_table_35 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pattern_table_36 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pattern_table_37 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pattern_table_38 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pattern_table_39 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pattern_table_40 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pattern_table_41 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pattern_table_42 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pattern_table_43 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pattern_table_44 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pattern_table_45 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pattern_table_46 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pattern_table_47 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pattern_table_48 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pattern_table_49 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pattern_table_50 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pattern_table_51 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pattern_table_52 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pattern_table_53 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pattern_table_54 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pattern_table_55 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pattern_table_56 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pattern_table_57 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pattern_table_58 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pattern_table_59 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pattern_table_60 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pattern_table_61 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pattern_table_62 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pattern_table_63 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pattern_table_64 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pattern_table_65 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pattern_table_66 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pattern_table_67 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pattern_table_68 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pattern_table_69 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pattern_table_70 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pattern_table_71 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pattern_table_72 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pattern_table_73 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pattern_table_74 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pattern_table_75 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pattern_table_76 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pattern_table_77 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pattern_table_78 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pattern_table_79 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pattern_table_80 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pattern_table_81 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pattern_table_82 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pattern_table_83 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pattern_table_84 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pattern_table_85 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pattern_table_86 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pattern_table_87 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pattern_table_88 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pattern_table_89 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pattern_table_90 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pattern_table_91 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pattern_table_92 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pattern_table_93 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pattern_table_94 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pattern_table_95 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pattern_table_96 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pattern_table_97 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pattern_table_98 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pattern_table_99 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pattern_table_100 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pattern_table_101 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pattern_table_102 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pattern_table_103 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pattern_table_104 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pattern_table_105 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pattern_table_106 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pattern_table_107 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pattern_table_108 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pattern_table_109 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pattern_table_110 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pattern_table_111 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pattern_table_112 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pattern_table_113 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pattern_table_114 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pattern_table_115 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pattern_table_116 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pattern_table_117 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pattern_table_118 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pattern_table_119 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pattern_table_120 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pattern_table_121 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pattern_table_122 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pattern_table_123 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pattern_table_124 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pattern_table_125 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pattern_table_126 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pattern_table_127 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pattern_table_128 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pattern_table_129 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pattern_table_130 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pattern_table_131 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pattern_table_132 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pattern_table_133 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pattern_table_134 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pattern_table_135 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pattern_table_136 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pattern_table_137 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pattern_table_138 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pattern_table_139 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pattern_table_140 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pattern_table_141 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pattern_table_142 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pattern_table_143 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pattern_table_144 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pattern_table_145 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pattern_table_146 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pattern_table_147 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pattern_table_148 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pattern_table_149 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pattern_table_150 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pattern_table_151 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pattern_table_152 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pattern_table_153 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pattern_table_154 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pattern_table_155 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pattern_table_156 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pattern_table_157 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pattern_table_158 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pattern_table_159 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pattern_table_160 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pattern_table_161 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pattern_table_162 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pattern_table_163 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pattern_table_164 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pattern_table_165 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pattern_table_166 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pattern_table_167 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pattern_table_168 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pattern_table_169 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pattern_table_170 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pattern_table_171 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pattern_table_172 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pattern_table_173 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pattern_table_174 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pattern_table_175 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pattern_table_176 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pattern_table_177 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pattern_table_178 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pattern_table_179 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pattern_table_180 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pattern_table_181 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pattern_table_182 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pattern_table_183 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pattern_table_184 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pattern_table_185 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pattern_table_186 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pattern_table_187 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pattern_table_188 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pattern_table_189 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pattern_table_190 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pattern_table_191 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pattern_table_192 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pattern_table_193 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pattern_table_194 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pattern_table_195 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pattern_table_196 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pattern_table_197 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pattern_table_198 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pattern_table_199 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pattern_table_200 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pattern_table_201 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pattern_table_202 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pattern_table_203 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pattern_table_204 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pattern_table_205 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pattern_table_206 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pattern_table_207 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pattern_table_208 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pattern_table_209 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pattern_table_210 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pattern_table_211 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pattern_table_212 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pattern_table_213 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pattern_table_214 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pattern_table_215 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pattern_table_216 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pattern_table_217 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pattern_table_218 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pattern_table_219 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pattern_table_220 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pattern_table_221 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pattern_table_222 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pattern_table_223 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pattern_table_224 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pattern_table_225 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pattern_table_226 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pattern_table_227 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pattern_table_228 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pattern_table_229 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pattern_table_230 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pattern_table_231 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pattern_table_232 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pattern_table_233 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pattern_table_234 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pattern_table_235 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pattern_table_236 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pattern_table_237 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pattern_table_238 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pattern_table_239 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pattern_table_240 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pattern_table_241 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pattern_table_242 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pattern_table_243 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pattern_table_244 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pattern_table_245 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pattern_table_246 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pattern_table_247 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pattern_table_248 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pattern_table_249 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pattern_table_250 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pattern_table_251 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pattern_table_252 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pattern_table_253 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pattern_table_254 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pattern_table_255 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  branch_target_buffer_0 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  branch_target_buffer_1 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  branch_target_buffer_2 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  branch_target_buffer_3 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  branch_target_buffer_4 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  branch_target_buffer_5 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  branch_target_buffer_6 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  branch_target_buffer_7 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  branch_target_buffer_8 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  branch_target_buffer_9 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  branch_target_buffer_10 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  branch_target_buffer_11 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  branch_target_buffer_12 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  branch_target_buffer_13 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  branch_target_buffer_14 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  branch_target_buffer_15 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  branch_target_buffer_16 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  branch_target_buffer_17 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  branch_target_buffer_18 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  branch_target_buffer_19 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  branch_target_buffer_20 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  branch_target_buffer_21 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  branch_target_buffer_22 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  branch_target_buffer_23 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  branch_target_buffer_24 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  branch_target_buffer_25 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  branch_target_buffer_26 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  branch_target_buffer_27 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  branch_target_buffer_28 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  branch_target_buffer_29 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  branch_target_buffer_30 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  branch_target_buffer_31 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  branch_target_buffer_32 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  branch_target_buffer_33 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  branch_target_buffer_34 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  branch_target_buffer_35 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  branch_target_buffer_36 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  branch_target_buffer_37 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  branch_target_buffer_38 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  branch_target_buffer_39 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  branch_target_buffer_40 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  branch_target_buffer_41 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  branch_target_buffer_42 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  branch_target_buffer_43 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  branch_target_buffer_44 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  branch_target_buffer_45 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  branch_target_buffer_46 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  branch_target_buffer_47 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  branch_target_buffer_48 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  branch_target_buffer_49 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  branch_target_buffer_50 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  branch_target_buffer_51 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  branch_target_buffer_52 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  branch_target_buffer_53 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  branch_target_buffer_54 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  branch_target_buffer_55 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  branch_target_buffer_56 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  branch_target_buffer_57 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  branch_target_buffer_58 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  branch_target_buffer_59 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  branch_target_buffer_60 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  branch_target_buffer_61 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  branch_target_buffer_62 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  branch_target_buffer_63 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  branch_target_buffer_64 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  branch_target_buffer_65 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  branch_target_buffer_66 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  branch_target_buffer_67 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  branch_target_buffer_68 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  branch_target_buffer_69 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  branch_target_buffer_70 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  branch_target_buffer_71 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  branch_target_buffer_72 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  branch_target_buffer_73 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  branch_target_buffer_74 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  branch_target_buffer_75 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  branch_target_buffer_76 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  branch_target_buffer_77 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  branch_target_buffer_78 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  branch_target_buffer_79 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  branch_target_buffer_80 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  branch_target_buffer_81 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  branch_target_buffer_82 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  branch_target_buffer_83 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  branch_target_buffer_84 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  branch_target_buffer_85 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  branch_target_buffer_86 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  branch_target_buffer_87 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  branch_target_buffer_88 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  branch_target_buffer_89 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  branch_target_buffer_90 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  branch_target_buffer_91 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  branch_target_buffer_92 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  branch_target_buffer_93 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  branch_target_buffer_94 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  branch_target_buffer_95 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  branch_target_buffer_96 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  branch_target_buffer_97 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  branch_target_buffer_98 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  branch_target_buffer_99 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  branch_target_buffer_100 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  branch_target_buffer_101 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  branch_target_buffer_102 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  branch_target_buffer_103 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  branch_target_buffer_104 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  branch_target_buffer_105 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  branch_target_buffer_106 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  branch_target_buffer_107 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  branch_target_buffer_108 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  branch_target_buffer_109 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  branch_target_buffer_110 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  branch_target_buffer_111 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  branch_target_buffer_112 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  branch_target_buffer_113 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  branch_target_buffer_114 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  branch_target_buffer_115 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  branch_target_buffer_116 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  branch_target_buffer_117 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  branch_target_buffer_118 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  branch_target_buffer_119 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  branch_target_buffer_120 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  branch_target_buffer_121 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  branch_target_buffer_122 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  branch_target_buffer_123 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  branch_target_buffer_124 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  branch_target_buffer_125 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  branch_target_buffer_126 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  branch_target_buffer_127 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  branch_target_buffer_128 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  branch_target_buffer_129 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  branch_target_buffer_130 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  branch_target_buffer_131 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  branch_target_buffer_132 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  branch_target_buffer_133 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  branch_target_buffer_134 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  branch_target_buffer_135 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  branch_target_buffer_136 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  branch_target_buffer_137 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  branch_target_buffer_138 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  branch_target_buffer_139 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  branch_target_buffer_140 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  branch_target_buffer_141 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  branch_target_buffer_142 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  branch_target_buffer_143 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  branch_target_buffer_144 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  branch_target_buffer_145 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  branch_target_buffer_146 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  branch_target_buffer_147 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  branch_target_buffer_148 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  branch_target_buffer_149 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  branch_target_buffer_150 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  branch_target_buffer_151 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  branch_target_buffer_152 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  branch_target_buffer_153 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  branch_target_buffer_154 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  branch_target_buffer_155 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  branch_target_buffer_156 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  branch_target_buffer_157 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  branch_target_buffer_158 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  branch_target_buffer_159 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  branch_target_buffer_160 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  branch_target_buffer_161 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  branch_target_buffer_162 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  branch_target_buffer_163 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  branch_target_buffer_164 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  branch_target_buffer_165 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  branch_target_buffer_166 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  branch_target_buffer_167 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  branch_target_buffer_168 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  branch_target_buffer_169 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  branch_target_buffer_170 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  branch_target_buffer_171 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  branch_target_buffer_172 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  branch_target_buffer_173 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  branch_target_buffer_174 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  branch_target_buffer_175 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  branch_target_buffer_176 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  branch_target_buffer_177 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  branch_target_buffer_178 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  branch_target_buffer_179 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  branch_target_buffer_180 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  branch_target_buffer_181 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  branch_target_buffer_182 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  branch_target_buffer_183 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  branch_target_buffer_184 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  branch_target_buffer_185 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  branch_target_buffer_186 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  branch_target_buffer_187 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  branch_target_buffer_188 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  branch_target_buffer_189 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  branch_target_buffer_190 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  branch_target_buffer_191 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  branch_target_buffer_192 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  branch_target_buffer_193 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  branch_target_buffer_194 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  branch_target_buffer_195 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  branch_target_buffer_196 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  branch_target_buffer_197 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  branch_target_buffer_198 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  branch_target_buffer_199 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  branch_target_buffer_200 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  branch_target_buffer_201 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  branch_target_buffer_202 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  branch_target_buffer_203 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  branch_target_buffer_204 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  branch_target_buffer_205 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  branch_target_buffer_206 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  branch_target_buffer_207 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  branch_target_buffer_208 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  branch_target_buffer_209 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  branch_target_buffer_210 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  branch_target_buffer_211 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  branch_target_buffer_212 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  branch_target_buffer_213 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  branch_target_buffer_214 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  branch_target_buffer_215 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  branch_target_buffer_216 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  branch_target_buffer_217 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  branch_target_buffer_218 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  branch_target_buffer_219 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  branch_target_buffer_220 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  branch_target_buffer_221 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  branch_target_buffer_222 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  branch_target_buffer_223 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  branch_target_buffer_224 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  branch_target_buffer_225 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  branch_target_buffer_226 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  branch_target_buffer_227 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  branch_target_buffer_228 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  branch_target_buffer_229 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  branch_target_buffer_230 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  branch_target_buffer_231 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  branch_target_buffer_232 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  branch_target_buffer_233 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  branch_target_buffer_234 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  branch_target_buffer_235 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  branch_target_buffer_236 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  branch_target_buffer_237 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  branch_target_buffer_238 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  branch_target_buffer_239 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  branch_target_buffer_240 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  branch_target_buffer_241 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  branch_target_buffer_242 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  branch_target_buffer_243 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  branch_target_buffer_244 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  branch_target_buffer_245 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  branch_target_buffer_246 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  branch_target_buffer_247 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  branch_target_buffer_248 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  branch_target_buffer_249 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  branch_target_buffer_250 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  branch_target_buffer_251 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  branch_target_buffer_252 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  branch_target_buffer_253 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  branch_target_buffer_254 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  branch_target_buffer_255 = _RAND_767[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ID(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_io_reg_pc,
  input  [31:0] io_in_if_io_inst,
  input         io_in_stall_io_stall_flag,
  input         io_in_stall_io_pred_miss_flag,
  input         io_in_mem_io_rd_wen,
  input  [4:0]  io_in_mem_io_rd_addr,
  input  [31:0] io_in_mem_io_rd_data,
  input         io_in_wb_io_rd_wen,
  input  [4:0]  io_in_wb_io_rd_addr,
  input  [31:0] io_in_wb_io_rd_data,
  output [31:0] io_out_op1_data,
  output [31:0] io_out_op2_data,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_csr_addr_default,
  output [4:0]  io_out_exe_fun,
  output        io_out_mem_wen,
  output        io_out_rd_wen,
  output [2:0]  io_out_rd_sel,
  output [2:0]  io_out_csr_cmd,
  output [31:0] io_out_rs2_data,
  output [31:0] io_out_imm_b_sext
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_x_0; // @[ID.scala 75:26]
  reg [31:0] reg_x_1; // @[ID.scala 75:26]
  reg [31:0] reg_x_2; // @[ID.scala 75:26]
  reg [31:0] reg_x_3; // @[ID.scala 75:26]
  reg [31:0] reg_x_4; // @[ID.scala 75:26]
  reg [31:0] reg_x_5; // @[ID.scala 75:26]
  reg [31:0] reg_x_6; // @[ID.scala 75:26]
  reg [31:0] reg_x_7; // @[ID.scala 75:26]
  reg [31:0] reg_x_8; // @[ID.scala 75:26]
  reg [31:0] reg_x_9; // @[ID.scala 75:26]
  reg [31:0] reg_x_10; // @[ID.scala 75:26]
  reg [31:0] reg_x_11; // @[ID.scala 75:26]
  reg [31:0] reg_x_12; // @[ID.scala 75:26]
  reg [31:0] reg_x_13; // @[ID.scala 75:26]
  reg [31:0] reg_x_14; // @[ID.scala 75:26]
  reg [31:0] reg_x_15; // @[ID.scala 75:26]
  reg [31:0] reg_x_16; // @[ID.scala 75:26]
  reg [31:0] reg_x_17; // @[ID.scala 75:26]
  reg [31:0] reg_x_18; // @[ID.scala 75:26]
  reg [31:0] reg_x_19; // @[ID.scala 75:26]
  reg [31:0] reg_x_20; // @[ID.scala 75:26]
  reg [31:0] reg_x_21; // @[ID.scala 75:26]
  reg [31:0] reg_x_22; // @[ID.scala 75:26]
  reg [31:0] reg_x_23; // @[ID.scala 75:26]
  reg [31:0] reg_x_24; // @[ID.scala 75:26]
  reg [31:0] reg_x_25; // @[ID.scala 75:26]
  reg [31:0] reg_x_26; // @[ID.scala 75:26]
  reg [31:0] reg_x_27; // @[ID.scala 75:26]
  reg [31:0] reg_x_28; // @[ID.scala 75:26]
  reg [31:0] reg_x_29; // @[ID.scala 75:26]
  reg [31:0] reg_x_30; // @[ID.scala 75:26]
  reg [31:0] reg_x_31; // @[ID.scala 75:26]
  wire [31:0] _inst_T = io_in_stall_io_stall_flag ? 32'h13 : io_in_if_io_inst; // @[Mux.scala 98:16]
  wire [31:0] inst = io_in_stall_io_pred_miss_flag ? 32'h13 : _inst_T; // @[Mux.scala 98:16]
  wire [4:0] rs1_addr = inst[19:15]; // @[ID.scala 95:24]
  wire [4:0] rs2_addr = inst[24:20]; // @[ID.scala 96:24]
  wire [4:0] rd_addr = inst[11:7]; // @[ID.scala 97:24]
  wire [11:0] csr_addr_default = inst[31:20]; // @[ID.scala 98:32]
  wire  _rs1_data_T = rs1_addr == 5'h0; // @[ID.scala 100:19]
  wire  _rs1_data_T_3 = rs1_addr == io_in_mem_io_rd_addr & io_in_mem_io_rd_wen; // @[ID.scala 101:37]
  wire  _rs1_data_T_6 = rs1_addr == io_in_wb_io_rd_addr & io_in_wb_io_rd_wen; // @[ID.scala 102:36]
  wire [31:0] _GEN_1 = 5'h1 == rs1_addr ? reg_x_1 : reg_x_0; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_2 = 5'h2 == rs1_addr ? reg_x_2 : _GEN_1; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_3 = 5'h3 == rs1_addr ? reg_x_3 : _GEN_2; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_4 = 5'h4 == rs1_addr ? reg_x_4 : _GEN_3; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_5 = 5'h5 == rs1_addr ? reg_x_5 : _GEN_4; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_6 = 5'h6 == rs1_addr ? reg_x_6 : _GEN_5; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_7 = 5'h7 == rs1_addr ? reg_x_7 : _GEN_6; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_8 = 5'h8 == rs1_addr ? reg_x_8 : _GEN_7; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_9 = 5'h9 == rs1_addr ? reg_x_9 : _GEN_8; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_10 = 5'ha == rs1_addr ? reg_x_10 : _GEN_9; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_11 = 5'hb == rs1_addr ? reg_x_11 : _GEN_10; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_12 = 5'hc == rs1_addr ? reg_x_12 : _GEN_11; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_13 = 5'hd == rs1_addr ? reg_x_13 : _GEN_12; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_14 = 5'he == rs1_addr ? reg_x_14 : _GEN_13; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_15 = 5'hf == rs1_addr ? reg_x_15 : _GEN_14; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_16 = 5'h10 == rs1_addr ? reg_x_16 : _GEN_15; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_17 = 5'h11 == rs1_addr ? reg_x_17 : _GEN_16; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_18 = 5'h12 == rs1_addr ? reg_x_18 : _GEN_17; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_19 = 5'h13 == rs1_addr ? reg_x_19 : _GEN_18; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_20 = 5'h14 == rs1_addr ? reg_x_20 : _GEN_19; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_21 = 5'h15 == rs1_addr ? reg_x_21 : _GEN_20; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_22 = 5'h16 == rs1_addr ? reg_x_22 : _GEN_21; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_23 = 5'h17 == rs1_addr ? reg_x_23 : _GEN_22; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_24 = 5'h18 == rs1_addr ? reg_x_24 : _GEN_23; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_25 = 5'h19 == rs1_addr ? reg_x_25 : _GEN_24; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_26 = 5'h1a == rs1_addr ? reg_x_26 : _GEN_25; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_27 = 5'h1b == rs1_addr ? reg_x_27 : _GEN_26; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_28 = 5'h1c == rs1_addr ? reg_x_28 : _GEN_27; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_29 = 5'h1d == rs1_addr ? reg_x_29 : _GEN_28; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_30 = 5'h1e == rs1_addr ? reg_x_30 : _GEN_29; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_31 = 5'h1f == rs1_addr ? reg_x_31 : _GEN_30; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _rs1_data_T_7 = _rs1_data_T_6 ? io_in_wb_io_rd_data : _GEN_31; // @[Mux.scala 98:16]
  wire [31:0] _rs1_data_T_8 = _rs1_data_T_3 ? io_in_mem_io_rd_data : _rs1_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] rs1_data = _rs1_data_T ? 32'h0 : _rs1_data_T_8; // @[Mux.scala 98:16]
  wire  _rs2_data_T = rs2_addr == 5'h0; // @[ID.scala 105:19]
  wire  _rs2_data_T_3 = rs2_addr == io_in_mem_io_rd_addr & io_in_mem_io_rd_wen; // @[ID.scala 106:37]
  wire  _rs2_data_T_6 = rs2_addr == io_in_wb_io_rd_addr & io_in_wb_io_rd_wen; // @[ID.scala 107:36]
  wire [31:0] _GEN_33 = 5'h1 == rs2_addr ? reg_x_1 : reg_x_0; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_34 = 5'h2 == rs2_addr ? reg_x_2 : _GEN_33; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_35 = 5'h3 == rs2_addr ? reg_x_3 : _GEN_34; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_36 = 5'h4 == rs2_addr ? reg_x_4 : _GEN_35; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_37 = 5'h5 == rs2_addr ? reg_x_5 : _GEN_36; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_38 = 5'h6 == rs2_addr ? reg_x_6 : _GEN_37; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_39 = 5'h7 == rs2_addr ? reg_x_7 : _GEN_38; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_40 = 5'h8 == rs2_addr ? reg_x_8 : _GEN_39; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_41 = 5'h9 == rs2_addr ? reg_x_9 : _GEN_40; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_42 = 5'ha == rs2_addr ? reg_x_10 : _GEN_41; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_43 = 5'hb == rs2_addr ? reg_x_11 : _GEN_42; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_44 = 5'hc == rs2_addr ? reg_x_12 : _GEN_43; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_45 = 5'hd == rs2_addr ? reg_x_13 : _GEN_44; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_46 = 5'he == rs2_addr ? reg_x_14 : _GEN_45; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_47 = 5'hf == rs2_addr ? reg_x_15 : _GEN_46; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_48 = 5'h10 == rs2_addr ? reg_x_16 : _GEN_47; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_49 = 5'h11 == rs2_addr ? reg_x_17 : _GEN_48; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_50 = 5'h12 == rs2_addr ? reg_x_18 : _GEN_49; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_51 = 5'h13 == rs2_addr ? reg_x_19 : _GEN_50; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_52 = 5'h14 == rs2_addr ? reg_x_20 : _GEN_51; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_53 = 5'h15 == rs2_addr ? reg_x_21 : _GEN_52; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_54 = 5'h16 == rs2_addr ? reg_x_22 : _GEN_53; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_55 = 5'h17 == rs2_addr ? reg_x_23 : _GEN_54; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_56 = 5'h18 == rs2_addr ? reg_x_24 : _GEN_55; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_57 = 5'h19 == rs2_addr ? reg_x_25 : _GEN_56; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_58 = 5'h1a == rs2_addr ? reg_x_26 : _GEN_57; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_59 = 5'h1b == rs2_addr ? reg_x_27 : _GEN_58; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_60 = 5'h1c == rs2_addr ? reg_x_28 : _GEN_59; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_61 = 5'h1d == rs2_addr ? reg_x_29 : _GEN_60; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_62 = 5'h1e == rs2_addr ? reg_x_30 : _GEN_61; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _GEN_63 = 5'h1f == rs2_addr ? reg_x_31 : _GEN_62; // @[Mux.scala 98:16 Mux.scala 98:16]
  wire [31:0] _rs2_data_T_7 = _rs2_data_T_6 ? io_in_wb_io_rd_data : _GEN_63; // @[Mux.scala 98:16]
  wire [31:0] _rs2_data_T_8 = _rs2_data_T_3 ? io_in_mem_io_rd_data : _rs2_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] rs2_data = _rs2_data_T ? 32'h0 : _rs2_data_T_8; // @[Mux.scala 98:16]
  wire [19:0] imm_i_sext_hi = csr_addr_default[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_i_sext = {imm_i_sext_hi,csr_addr_default}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi = inst[31:25]; // @[ID.scala 111:31]
  wire [11:0] imm_s = {imm_s_hi,rd_addr}; // @[Cat.scala 30:58]
  wire [19:0] imm_s_sext_hi = imm_s[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_s_sext = {imm_s_sext_hi,imm_s_hi,rd_addr}; // @[Cat.scala 30:58]
  wire  imm_b_hi_hi = inst[31]; // @[ID.scala 113:31]
  wire  imm_b_hi_lo = inst[7]; // @[ID.scala 113:41]
  wire [5:0] imm_b_lo_hi = inst[30:25]; // @[ID.scala 113:50]
  wire [3:0] imm_b_lo_lo = inst[11:8]; // @[ID.scala 113:64]
  wire [11:0] imm_b = {imm_b_hi_hi,imm_b_hi_lo,imm_b_lo_hi,imm_b_lo_lo}; // @[Cat.scala 30:58]
  wire [18:0] imm_b_sext_hi_hi = imm_b[11] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [30:0] imm_b_sext_hi = {imm_b_sext_hi_hi,imm_b_hi_hi,imm_b_hi_lo,imm_b_lo_hi,imm_b_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] imm_j_hi_lo = inst[19:12]; // @[ID.scala 115:41]
  wire  imm_j_lo_hi = inst[20]; // @[ID.scala 115:55]
  wire [9:0] imm_j_lo_lo = inst[30:21]; // @[ID.scala 115:65]
  wire [19:0] imm_j = {imm_b_hi_hi,imm_j_hi_lo,imm_j_lo_hi,imm_j_lo_lo}; // @[Cat.scala 30:58]
  wire [10:0] imm_j_sext_hi_hi = imm_j[19] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_j_sext = {imm_j_sext_hi_hi,imm_b_hi_hi,imm_j_hi_lo,imm_j_lo_hi,imm_j_lo_lo,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] imm_u = inst[31:12]; // @[ID.scala 117:27]
  wire [31:0] imm_u_shifted = {imm_u,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_z_uext = {27'h0,rs1_addr}; // @[Cat.scala 30:58]
  wire [31:0] _inst_type_T = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_1 = 32'h2003 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_3 = 32'h2023 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_4 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_5 = 32'h33 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_7 = 32'h13 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_9 = 32'h40000033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_11 = 32'h7033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_13 = 32'h6033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_15 = 32'h4033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_17 = 32'h7013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_19 = 32'h6013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_21 = 32'h4013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_23 = 32'h1033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_25 = 32'h5033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_27 = 32'h40005033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_29 = 32'h1013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_31 = 32'h5013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_33 = 32'h40005013 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_35 = 32'h2033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_37 = 32'h3033 == _inst_type_T_4; // @[Lookup.scala 31:38]
  wire  _inst_type_T_39 = 32'h2013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_41 = 32'h3013 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_43 = 32'h63 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_45 = 32'h1063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_47 = 32'h5063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_49 = 32'h7063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_51 = 32'h4063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_53 = 32'h6063 == _inst_type_T; // @[Lookup.scala 31:38]
  wire [31:0] _inst_type_T_54 = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _inst_type_T_55 = 32'h6f == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_57 = 32'h67 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_59 = 32'h37 == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_61 = 32'h17 == _inst_type_T_54; // @[Lookup.scala 31:38]
  wire  _inst_type_T_63 = 32'h1073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_65 = 32'h5073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_67 = 32'h2073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_69 = 32'h6073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_71 = 32'h3073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_73 = 32'h7073 == _inst_type_T; // @[Lookup.scala 31:38]
  wire  _inst_type_T_75 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire [4:0] _inst_type_T_77 = _inst_type_T_73 ? 5'h12 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_78 = _inst_type_T_71 ? 5'h12 : _inst_type_T_77; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_79 = _inst_type_T_69 ? 5'h12 : _inst_type_T_78; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_80 = _inst_type_T_67 ? 5'h12 : _inst_type_T_79; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_81 = _inst_type_T_65 ? 5'h12 : _inst_type_T_80; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_82 = _inst_type_T_63 ? 5'h12 : _inst_type_T_81; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_83 = _inst_type_T_61 ? 5'h1 : _inst_type_T_82; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_84 = _inst_type_T_59 ? 5'h1 : _inst_type_T_83; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_85 = _inst_type_T_57 ? 5'h11 : _inst_type_T_84; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_86 = _inst_type_T_55 ? 5'h1 : _inst_type_T_85; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_87 = _inst_type_T_53 ? 5'hf : _inst_type_T_86; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_88 = _inst_type_T_51 ? 5'hd : _inst_type_T_87; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_89 = _inst_type_T_49 ? 5'h10 : _inst_type_T_88; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_90 = _inst_type_T_47 ? 5'he : _inst_type_T_89; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_91 = _inst_type_T_45 ? 5'hc : _inst_type_T_90; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_92 = _inst_type_T_43 ? 5'hb : _inst_type_T_91; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_93 = _inst_type_T_41 ? 5'ha : _inst_type_T_92; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_94 = _inst_type_T_39 ? 5'h9 : _inst_type_T_93; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_95 = _inst_type_T_37 ? 5'ha : _inst_type_T_94; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_96 = _inst_type_T_35 ? 5'h9 : _inst_type_T_95; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_97 = _inst_type_T_33 ? 5'h8 : _inst_type_T_96; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_98 = _inst_type_T_31 ? 5'h7 : _inst_type_T_97; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_99 = _inst_type_T_29 ? 5'h6 : _inst_type_T_98; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_100 = _inst_type_T_27 ? 5'h8 : _inst_type_T_99; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_101 = _inst_type_T_25 ? 5'h7 : _inst_type_T_100; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_102 = _inst_type_T_23 ? 5'h6 : _inst_type_T_101; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_103 = _inst_type_T_21 ? 5'h5 : _inst_type_T_102; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_104 = _inst_type_T_19 ? 5'h4 : _inst_type_T_103; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_105 = _inst_type_T_17 ? 5'h3 : _inst_type_T_104; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_106 = _inst_type_T_15 ? 5'h5 : _inst_type_T_105; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_107 = _inst_type_T_13 ? 5'h4 : _inst_type_T_106; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_108 = _inst_type_T_11 ? 5'h3 : _inst_type_T_107; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_109 = _inst_type_T_9 ? 5'h2 : _inst_type_T_108; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_110 = _inst_type_T_7 ? 5'h1 : _inst_type_T_109; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_111 = _inst_type_T_5 ? 5'h1 : _inst_type_T_110; // @[Lookup.scala 33:37]
  wire [4:0] _inst_type_T_112 = _inst_type_T_3 ? 5'h1 : _inst_type_T_111; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_113 = _inst_type_T_75 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_114 = _inst_type_T_73 ? 2'h3 : _inst_type_T_113; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_115 = _inst_type_T_71 ? 2'h0 : _inst_type_T_114; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_116 = _inst_type_T_69 ? 2'h3 : _inst_type_T_115; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_117 = _inst_type_T_67 ? 2'h0 : _inst_type_T_116; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_118 = _inst_type_T_65 ? 2'h3 : _inst_type_T_117; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_119 = _inst_type_T_63 ? 2'h0 : _inst_type_T_118; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_120 = _inst_type_T_61 ? 2'h1 : _inst_type_T_119; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_121 = _inst_type_T_59 ? 2'h2 : _inst_type_T_120; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_122 = _inst_type_T_57 ? 2'h0 : _inst_type_T_121; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_123 = _inst_type_T_55 ? 2'h1 : _inst_type_T_122; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_124 = _inst_type_T_53 ? 2'h0 : _inst_type_T_123; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_125 = _inst_type_T_51 ? 2'h0 : _inst_type_T_124; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_126 = _inst_type_T_49 ? 2'h0 : _inst_type_T_125; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_127 = _inst_type_T_47 ? 2'h0 : _inst_type_T_126; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_128 = _inst_type_T_45 ? 2'h0 : _inst_type_T_127; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_129 = _inst_type_T_43 ? 2'h0 : _inst_type_T_128; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_130 = _inst_type_T_41 ? 2'h0 : _inst_type_T_129; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_131 = _inst_type_T_39 ? 2'h0 : _inst_type_T_130; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_132 = _inst_type_T_37 ? 2'h0 : _inst_type_T_131; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_133 = _inst_type_T_35 ? 2'h0 : _inst_type_T_132; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_134 = _inst_type_T_33 ? 2'h0 : _inst_type_T_133; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_135 = _inst_type_T_31 ? 2'h0 : _inst_type_T_134; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_136 = _inst_type_T_29 ? 2'h0 : _inst_type_T_135; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_137 = _inst_type_T_27 ? 2'h0 : _inst_type_T_136; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_138 = _inst_type_T_25 ? 2'h0 : _inst_type_T_137; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_139 = _inst_type_T_23 ? 2'h0 : _inst_type_T_138; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_140 = _inst_type_T_21 ? 2'h0 : _inst_type_T_139; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_141 = _inst_type_T_19 ? 2'h0 : _inst_type_T_140; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_142 = _inst_type_T_17 ? 2'h0 : _inst_type_T_141; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_143 = _inst_type_T_15 ? 2'h0 : _inst_type_T_142; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_144 = _inst_type_T_13 ? 2'h0 : _inst_type_T_143; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_145 = _inst_type_T_11 ? 2'h0 : _inst_type_T_144; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_146 = _inst_type_T_9 ? 2'h0 : _inst_type_T_145; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_147 = _inst_type_T_7 ? 2'h0 : _inst_type_T_146; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_148 = _inst_type_T_5 ? 2'h0 : _inst_type_T_147; // @[Lookup.scala 33:37]
  wire [1:0] _inst_type_T_149 = _inst_type_T_3 ? 2'h0 : _inst_type_T_148; // @[Lookup.scala 33:37]
  wire [1:0] inst_type_1 = _inst_type_T_1 ? 2'h0 : _inst_type_T_149; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_150 = _inst_type_T_75 ? 3'h0 : 3'h1; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_151 = _inst_type_T_73 ? 3'h0 : _inst_type_T_150; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_152 = _inst_type_T_71 ? 3'h0 : _inst_type_T_151; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_153 = _inst_type_T_69 ? 3'h0 : _inst_type_T_152; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_154 = _inst_type_T_67 ? 3'h0 : _inst_type_T_153; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_155 = _inst_type_T_65 ? 3'h0 : _inst_type_T_154; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_156 = _inst_type_T_63 ? 3'h0 : _inst_type_T_155; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_157 = _inst_type_T_61 ? 3'h5 : _inst_type_T_156; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_158 = _inst_type_T_59 ? 3'h5 : _inst_type_T_157; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_159 = _inst_type_T_57 ? 3'h2 : _inst_type_T_158; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_160 = _inst_type_T_55 ? 3'h4 : _inst_type_T_159; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_161 = _inst_type_T_53 ? 3'h1 : _inst_type_T_160; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_162 = _inst_type_T_51 ? 3'h1 : _inst_type_T_161; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_163 = _inst_type_T_49 ? 3'h1 : _inst_type_T_162; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_164 = _inst_type_T_47 ? 3'h1 : _inst_type_T_163; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_165 = _inst_type_T_45 ? 3'h1 : _inst_type_T_164; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_166 = _inst_type_T_43 ? 3'h1 : _inst_type_T_165; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_167 = _inst_type_T_41 ? 3'h2 : _inst_type_T_166; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_168 = _inst_type_T_39 ? 3'h2 : _inst_type_T_167; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_169 = _inst_type_T_37 ? 3'h1 : _inst_type_T_168; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_170 = _inst_type_T_35 ? 3'h1 : _inst_type_T_169; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_171 = _inst_type_T_33 ? 3'h2 : _inst_type_T_170; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_172 = _inst_type_T_31 ? 3'h2 : _inst_type_T_171; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_173 = _inst_type_T_29 ? 3'h2 : _inst_type_T_172; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_174 = _inst_type_T_27 ? 3'h1 : _inst_type_T_173; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_175 = _inst_type_T_25 ? 3'h1 : _inst_type_T_174; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_176 = _inst_type_T_23 ? 3'h1 : _inst_type_T_175; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_177 = _inst_type_T_21 ? 3'h2 : _inst_type_T_176; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_178 = _inst_type_T_19 ? 3'h2 : _inst_type_T_177; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_179 = _inst_type_T_17 ? 3'h2 : _inst_type_T_178; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_180 = _inst_type_T_15 ? 3'h1 : _inst_type_T_179; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_181 = _inst_type_T_13 ? 3'h1 : _inst_type_T_180; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_182 = _inst_type_T_11 ? 3'h1 : _inst_type_T_181; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_183 = _inst_type_T_9 ? 3'h1 : _inst_type_T_182; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_184 = _inst_type_T_7 ? 3'h2 : _inst_type_T_183; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_185 = _inst_type_T_5 ? 3'h1 : _inst_type_T_184; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_186 = _inst_type_T_3 ? 3'h3 : _inst_type_T_185; // @[Lookup.scala 33:37]
  wire [2:0] inst_type_2 = _inst_type_T_1 ? 3'h2 : _inst_type_T_186; // @[Lookup.scala 33:37]
  wire  _inst_type_T_235 = _inst_type_T_53 ? 1'h0 : _inst_type_T_55 | (_inst_type_T_57 | (_inst_type_T_59 | (
    _inst_type_T_61 | (_inst_type_T_63 | (_inst_type_T_65 | (_inst_type_T_67 | (_inst_type_T_69 | (_inst_type_T_71 |
    _inst_type_T_73)))))))); // @[Lookup.scala 33:37]
  wire  _inst_type_T_236 = _inst_type_T_51 ? 1'h0 : _inst_type_T_235; // @[Lookup.scala 33:37]
  wire  _inst_type_T_237 = _inst_type_T_49 ? 1'h0 : _inst_type_T_236; // @[Lookup.scala 33:37]
  wire  _inst_type_T_238 = _inst_type_T_47 ? 1'h0 : _inst_type_T_237; // @[Lookup.scala 33:37]
  wire  _inst_type_T_239 = _inst_type_T_45 ? 1'h0 : _inst_type_T_238; // @[Lookup.scala 33:37]
  wire  _inst_type_T_240 = _inst_type_T_43 ? 1'h0 : _inst_type_T_239; // @[Lookup.scala 33:37]
  wire  _inst_type_T_260 = _inst_type_T_3 ? 1'h0 : _inst_type_T_5 | (_inst_type_T_7 | (_inst_type_T_9 | (_inst_type_T_11
     | (_inst_type_T_13 | (_inst_type_T_15 | (_inst_type_T_17 | (_inst_type_T_19 | (_inst_type_T_21 | (_inst_type_T_23
     | (_inst_type_T_25 | (_inst_type_T_27 | (_inst_type_T_29 | (_inst_type_T_31 | (_inst_type_T_33 | (_inst_type_T_35
     | (_inst_type_T_37 | (_inst_type_T_39 | (_inst_type_T_41 | _inst_type_T_240)))))))))))))))))); // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_262 = _inst_type_T_73 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_263 = _inst_type_T_71 ? 3'h3 : _inst_type_T_262; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_264 = _inst_type_T_69 ? 3'h3 : _inst_type_T_263; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_265 = _inst_type_T_67 ? 3'h3 : _inst_type_T_264; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_266 = _inst_type_T_65 ? 3'h3 : _inst_type_T_265; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_267 = _inst_type_T_63 ? 3'h3 : _inst_type_T_266; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_268 = _inst_type_T_61 ? 3'h0 : _inst_type_T_267; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_269 = _inst_type_T_59 ? 3'h0 : _inst_type_T_268; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_270 = _inst_type_T_57 ? 3'h2 : _inst_type_T_269; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_271 = _inst_type_T_55 ? 3'h2 : _inst_type_T_270; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_272 = _inst_type_T_53 ? 3'h0 : _inst_type_T_271; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_273 = _inst_type_T_51 ? 3'h0 : _inst_type_T_272; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_274 = _inst_type_T_49 ? 3'h0 : _inst_type_T_273; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_275 = _inst_type_T_47 ? 3'h0 : _inst_type_T_274; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_276 = _inst_type_T_45 ? 3'h0 : _inst_type_T_275; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_277 = _inst_type_T_43 ? 3'h0 : _inst_type_T_276; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_278 = _inst_type_T_41 ? 3'h0 : _inst_type_T_277; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_279 = _inst_type_T_39 ? 3'h0 : _inst_type_T_278; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_280 = _inst_type_T_37 ? 3'h0 : _inst_type_T_279; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_281 = _inst_type_T_35 ? 3'h0 : _inst_type_T_280; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_282 = _inst_type_T_33 ? 3'h0 : _inst_type_T_281; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_283 = _inst_type_T_31 ? 3'h0 : _inst_type_T_282; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_284 = _inst_type_T_29 ? 3'h0 : _inst_type_T_283; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_285 = _inst_type_T_27 ? 3'h0 : _inst_type_T_284; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_286 = _inst_type_T_25 ? 3'h0 : _inst_type_T_285; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_287 = _inst_type_T_23 ? 3'h0 : _inst_type_T_286; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_288 = _inst_type_T_21 ? 3'h0 : _inst_type_T_287; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_289 = _inst_type_T_19 ? 3'h0 : _inst_type_T_288; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_290 = _inst_type_T_17 ? 3'h0 : _inst_type_T_289; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_291 = _inst_type_T_15 ? 3'h0 : _inst_type_T_290; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_292 = _inst_type_T_13 ? 3'h0 : _inst_type_T_291; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_293 = _inst_type_T_11 ? 3'h0 : _inst_type_T_292; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_294 = _inst_type_T_9 ? 3'h0 : _inst_type_T_293; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_295 = _inst_type_T_7 ? 3'h0 : _inst_type_T_294; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_296 = _inst_type_T_5 ? 3'h0 : _inst_type_T_295; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_297 = _inst_type_T_3 ? 3'h0 : _inst_type_T_296; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_298 = _inst_type_T_75 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_299 = _inst_type_T_73 ? 3'h3 : _inst_type_T_298; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_300 = _inst_type_T_71 ? 3'h3 : _inst_type_T_299; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_301 = _inst_type_T_69 ? 3'h2 : _inst_type_T_300; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_302 = _inst_type_T_67 ? 3'h2 : _inst_type_T_301; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_303 = _inst_type_T_65 ? 3'h1 : _inst_type_T_302; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_304 = _inst_type_T_63 ? 3'h1 : _inst_type_T_303; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_305 = _inst_type_T_61 ? 3'h0 : _inst_type_T_304; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_306 = _inst_type_T_59 ? 3'h0 : _inst_type_T_305; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_307 = _inst_type_T_57 ? 3'h0 : _inst_type_T_306; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_308 = _inst_type_T_55 ? 3'h0 : _inst_type_T_307; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_309 = _inst_type_T_53 ? 3'h0 : _inst_type_T_308; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_310 = _inst_type_T_51 ? 3'h0 : _inst_type_T_309; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_311 = _inst_type_T_49 ? 3'h0 : _inst_type_T_310; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_312 = _inst_type_T_47 ? 3'h0 : _inst_type_T_311; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_313 = _inst_type_T_45 ? 3'h0 : _inst_type_T_312; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_314 = _inst_type_T_43 ? 3'h0 : _inst_type_T_313; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_315 = _inst_type_T_41 ? 3'h0 : _inst_type_T_314; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_316 = _inst_type_T_39 ? 3'h0 : _inst_type_T_315; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_317 = _inst_type_T_37 ? 3'h0 : _inst_type_T_316; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_318 = _inst_type_T_35 ? 3'h0 : _inst_type_T_317; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_319 = _inst_type_T_33 ? 3'h0 : _inst_type_T_318; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_320 = _inst_type_T_31 ? 3'h0 : _inst_type_T_319; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_321 = _inst_type_T_29 ? 3'h0 : _inst_type_T_320; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_322 = _inst_type_T_27 ? 3'h0 : _inst_type_T_321; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_323 = _inst_type_T_25 ? 3'h0 : _inst_type_T_322; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_324 = _inst_type_T_23 ? 3'h0 : _inst_type_T_323; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_325 = _inst_type_T_21 ? 3'h0 : _inst_type_T_324; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_326 = _inst_type_T_19 ? 3'h0 : _inst_type_T_325; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_327 = _inst_type_T_17 ? 3'h0 : _inst_type_T_326; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_328 = _inst_type_T_15 ? 3'h0 : _inst_type_T_327; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_329 = _inst_type_T_13 ? 3'h0 : _inst_type_T_328; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_330 = _inst_type_T_11 ? 3'h0 : _inst_type_T_329; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_331 = _inst_type_T_9 ? 3'h0 : _inst_type_T_330; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_332 = _inst_type_T_7 ? 3'h0 : _inst_type_T_331; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_333 = _inst_type_T_5 ? 3'h0 : _inst_type_T_332; // @[Lookup.scala 33:37]
  wire [2:0] _inst_type_T_334 = _inst_type_T_3 ? 3'h0 : _inst_type_T_333; // @[Lookup.scala 33:37]
  wire  _op1_data_T = inst_type_1 == 2'h0; // @[ID.scala 168:18]
  wire  _op1_data_T_1 = inst_type_1 == 2'h1; // @[ID.scala 169:18]
  wire  _op1_data_T_2 = inst_type_1 == 2'h3; // @[ID.scala 170:18]
  wire [31:0] _op1_data_T_3 = _op1_data_T_2 ? imm_z_uext : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _op1_data_T_4 = _op1_data_T_1 ? io_in_if_io_reg_pc : _op1_data_T_3; // @[Mux.scala 98:16]
  wire [31:0] op1_data = _op1_data_T ? rs1_data : _op1_data_T_4; // @[Mux.scala 98:16]
  wire  _op2_data_T = inst_type_2 == 3'h1; // @[ID.scala 174:18]
  wire  _op2_data_T_1 = inst_type_2 == 3'h2; // @[ID.scala 175:18]
  wire  _op2_data_T_2 = inst_type_2 == 3'h3; // @[ID.scala 176:18]
  wire  _op2_data_T_3 = inst_type_2 == 3'h4; // @[ID.scala 177:18]
  wire  _op2_data_T_4 = inst_type_2 == 3'h5; // @[ID.scala 178:18]
  wire [31:0] _op2_data_T_5 = _op2_data_T_4 ? imm_u_shifted : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_6 = _op2_data_T_3 ? imm_j_sext : _op2_data_T_5; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_7 = _op2_data_T_2 ? imm_s_sext : _op2_data_T_6; // @[Mux.scala 98:16]
  wire [31:0] _op2_data_T_8 = _op2_data_T_1 ? imm_i_sext : _op2_data_T_7; // @[Mux.scala 98:16]
  wire [31:0] op2_data = _op2_data_T ? rs2_data : _op2_data_T_8; // @[Mux.scala 98:16]
  wire [31:0] _GEN_128 = {{27'd0}, io_in_wb_io_rd_addr}; // @[ID.scala 182:45]
  wire  _T_4 = ~reset; // @[ID.scala 202:11]
  assign io_out_op1_data = _op1_data_T ? rs1_data : _op1_data_T_4; // @[Mux.scala 98:16]
  assign io_out_op2_data = _op2_data_T ? rs2_data : _op2_data_T_8; // @[Mux.scala 98:16]
  assign io_out_rd_addr = inst[11:7]; // @[ID.scala 97:24]
  assign io_out_csr_addr_default = {{20'd0}, csr_addr_default}; // @[ID.scala 98:32]
  assign io_out_exe_fun = _inst_type_T_1 ? 5'h1 : _inst_type_T_112; // @[Lookup.scala 33:37]
  assign io_out_mem_wen = _inst_type_T_1 ? 1'h0 : _inst_type_T_3; // @[Lookup.scala 33:37]
  assign io_out_rd_wen = _inst_type_T_1 | _inst_type_T_260; // @[Lookup.scala 33:37]
  assign io_out_rd_sel = _inst_type_T_1 ? 3'h1 : _inst_type_T_297; // @[Lookup.scala 33:37]
  assign io_out_csr_cmd = _inst_type_T_1 ? 3'h0 : _inst_type_T_334; // @[Lookup.scala 33:37]
  assign io_out_rs2_data = _rs2_data_T ? 32'h0 : _rs2_data_T_8; // @[Mux.scala 98:16]
  assign io_out_imm_b_sext = {imm_b_sext_hi,1'h0}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[ID.scala 75:26]
      reg_x_0 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h0 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_0 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_1 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_1 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_2 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h2 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_2 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_3 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h3 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_3 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_4 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h4 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_4 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_5 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h5 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_5 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_6 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h6 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_6 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_7 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h7 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_7 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_8 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h8 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_8 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_9 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h9 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_9 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_10 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'ha == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_10 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_11 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hb == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_11 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_12 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hc == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_12 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_13 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hd == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_13 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_14 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'he == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_14 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_15 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'hf == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_15 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_16 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h10 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_16 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_17 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h11 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_17 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_18 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h12 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_18 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_19 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h13 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_19 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_20 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h14 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_20 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_21 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h15 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_21 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_22 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h16 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_22 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_23 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h17 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_23 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_24 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h18 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_24 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_25 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h19 == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_25 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_26 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1a == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_26 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_27 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1b == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_27 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_28 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1c == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_28 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_29 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1d == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_29 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_30 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1e == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_30 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    if (reset) begin // @[ID.scala 75:26]
      reg_x_31 <= 32'h0; // @[ID.scala 75:26]
    end else if (io_in_wb_io_rd_wen & _GEN_128 != 32'h0) begin // @[ID.scala 182:65]
      if (5'h1f == io_in_wb_io_rd_addr) begin // @[ID.scala 183:27]
        reg_x_31 <= io_in_wb_io_rd_data; // @[ID.scala 183:27]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------ID------------\n"); // @[ID.scala 202:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"rs1_addr: %d\n",rs1_addr); // @[ID.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"rs2_addr: %d\n",rs2_addr); // @[ID.scala 204:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"op1_data: 0x%x\n",op1_data); // @[ID.scala 205:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"op2_data: 0x%x\n",op2_data); // @[ID.scala 206:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"stall_flag: %d\n",io_in_stall_io_stall_flag); // @[ID.scala 207:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_x_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_x_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_x_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_x_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_x_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_x_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_x_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_x_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_x_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_x_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_x_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_x_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_x_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_x_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_x_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_x_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_x_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_x_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_x_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_x_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_x_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_x_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_x_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_x_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_x_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_x_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_x_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_x_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_x_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_x_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_x_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_x_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Stall(
  input  [31:0] io_in_if_io_reg_pc,
  input  [31:0] io_in_if_io_inst,
  input  [31:0] io_in_if_io_ex_io_alu_io_alu_out,
  input         io_in_if_io_ex_io_alu_io_jump_flag,
  input         io_in_if_io_ex_io_br_io_br_flag,
  input  [31:0] io_in_if_io_ex_io_br_io_br_target,
  input  [4:0]  io_in_id_reg_io_rd_addr,
  input         io_in_id_reg_io_rd_wen,
  output        io_out_stall_flag,
  output        io_out_pred_miss_flag
);
  wire [4:0] rs1_addr_default = io_in_if_io_inst[19:15]; // @[Stall.scala 42:43]
  wire [4:0] rs2_addr_default = io_in_if_io_inst[24:20]; // @[Stall.scala 43:43]
  wire  rs1_data_hazard = io_in_id_reg_io_rd_wen & rs1_addr_default != 5'h0 & rs1_addr_default ==
    io_in_id_reg_io_rd_addr; // @[Stall.scala 44:84]
  wire  rs2_data_hazard = io_in_id_reg_io_rd_wen & rs2_addr_default != 5'h0 & rs2_addr_default ==
    io_in_id_reg_io_rd_addr; // @[Stall.scala 45:84]
  assign io_out_stall_flag = rs1_data_hazard | rs2_data_hazard; // @[Stall.scala 46:48]
  assign io_out_pred_miss_flag = io_in_if_io_ex_io_alu_io_jump_flag & io_in_if_io_reg_pc !=
    io_in_if_io_ex_io_alu_io_alu_out | io_in_if_io_ex_io_br_io_br_flag & io_in_if_io_reg_pc !=
    io_in_if_io_ex_io_br_io_br_target; // @[Stall.scala 47:71]
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_in_id_io_op1_data,
  input  [31:0] io_in_id_io_op2_data,
  input  [4:0]  io_in_id_io_exe_fun,
  input  [2:0]  io_in_id_io_rd_sel,
  output [31:0] io_out_alu_out,
  output        io_out_jump_flag
);
  wire  _alu_out_T = io_in_id_io_exe_fun == 5'h1; // @[ALU.scala 38:18]
  wire [31:0] _alu_out_T_2 = io_in_id_io_op1_data + io_in_id_io_op2_data; // @[ALU.scala 38:46]
  wire  _alu_out_T_3 = io_in_id_io_exe_fun == 5'h2; // @[ALU.scala 39:18]
  wire [31:0] _alu_out_T_5 = io_in_id_io_op1_data - io_in_id_io_op2_data; // @[ALU.scala 39:46]
  wire  _alu_out_T_6 = io_in_id_io_exe_fun == 5'h3; // @[ALU.scala 40:18]
  wire [31:0] _alu_out_T_7 = io_in_id_io_op1_data & io_in_id_io_op2_data; // @[ALU.scala 40:46]
  wire  _alu_out_T_8 = io_in_id_io_exe_fun == 5'h4; // @[ALU.scala 41:18]
  wire [31:0] _alu_out_T_9 = io_in_id_io_op1_data | io_in_id_io_op2_data; // @[ALU.scala 41:46]
  wire  _alu_out_T_10 = io_in_id_io_exe_fun == 5'h5; // @[ALU.scala 42:18]
  wire [31:0] _alu_out_T_11 = io_in_id_io_op1_data ^ io_in_id_io_op2_data; // @[ALU.scala 42:46]
  wire  _alu_out_T_12 = io_in_id_io_exe_fun == 5'h6; // @[ALU.scala 43:18]
  wire [62:0] _GEN_0 = {{31'd0}, io_in_id_io_op1_data}; // @[ALU.scala 43:46]
  wire [62:0] _alu_out_T_14 = _GEN_0 << io_in_id_io_op2_data[4:0]; // @[ALU.scala 43:46]
  wire  _alu_out_T_16 = io_in_id_io_exe_fun == 5'h7; // @[ALU.scala 44:18]
  wire [31:0] _alu_out_T_18 = io_in_id_io_op1_data >> io_in_id_io_op2_data[4:0]; // @[ALU.scala 44:46]
  wire  _alu_out_T_19 = io_in_id_io_exe_fun == 5'h8; // @[ALU.scala 45:18]
  wire [31:0] _alu_out_T_23 = $signed(io_in_id_io_op1_data) >>> io_in_id_io_op2_data[4:0]; // @[ALU.scala 45:80]
  wire  _alu_out_T_24 = io_in_id_io_exe_fun == 5'h9; // @[ALU.scala 46:18]
  wire  _alu_out_T_27 = $signed(io_in_id_io_op1_data) < $signed(io_in_id_io_op2_data); // @[ALU.scala 46:55]
  wire  _alu_out_T_28 = io_in_id_io_exe_fun == 5'ha; // @[ALU.scala 47:18]
  wire  _alu_out_T_29 = io_in_id_io_op1_data < io_in_id_io_op2_data; // @[ALU.scala 47:46]
  wire  _alu_out_T_30 = io_in_id_io_exe_fun == 5'h11; // @[ALU.scala 48:18]
  wire [31:0] _alu_out_T_34 = _alu_out_T_2 & 32'hfffffffe; // @[ALU.scala 48:59]
  wire  _alu_out_T_35 = io_in_id_io_exe_fun == 5'h12; // @[ALU.scala 49:18]
  wire [31:0] _alu_out_T_36 = _alu_out_T_35 ? io_in_id_io_op1_data : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_37 = _alu_out_T_30 ? _alu_out_T_34 : _alu_out_T_36; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_38 = _alu_out_T_28 ? {{31'd0}, _alu_out_T_29} : _alu_out_T_37; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_39 = _alu_out_T_24 ? {{31'd0}, _alu_out_T_27} : _alu_out_T_38; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_40 = _alu_out_T_19 ? _alu_out_T_23 : _alu_out_T_39; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_41 = _alu_out_T_16 ? _alu_out_T_18 : _alu_out_T_40; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_42 = _alu_out_T_12 ? _alu_out_T_14[31:0] : _alu_out_T_41; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_43 = _alu_out_T_10 ? _alu_out_T_11 : _alu_out_T_42; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_44 = _alu_out_T_8 ? _alu_out_T_9 : _alu_out_T_43; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_45 = _alu_out_T_6 ? _alu_out_T_7 : _alu_out_T_44; // @[Mux.scala 98:16]
  wire [31:0] _alu_out_T_46 = _alu_out_T_3 ? _alu_out_T_5 : _alu_out_T_45; // @[Mux.scala 98:16]
  wire [31:0] alu_out = _alu_out_T ? _alu_out_T_2 : _alu_out_T_46; // @[Mux.scala 98:16]
  wire  jump_flag = io_in_id_io_rd_sel == 3'h2; // @[ALU.scala 52:29]
  wire  _T_1 = ~reset; // @[ALU.scala 59:11]
  assign io_out_alu_out = _alu_out_T ? _alu_out_T_2 : _alu_out_T_46; // @[Mux.scala 98:16]
  assign io_out_jump_flag = io_in_id_io_rd_sel == 3'h2; // @[ALU.scala 52:29]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------EX------------\n"); // @[ALU.scala 59:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"alu_out: 0x%x\n",alu_out); // @[ALU.scala 60:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"jump_flg: %d\n",jump_flag); // @[ALU.scala 61:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [31:0] io_in_id_io_op1_data,
  input  [31:0] io_in_id_io_csr_addr_default,
  input  [2:0]  io_in_id_io_csr_cmd,
  output [31:0] io_out_csr_rdata,
  output [31:0] io_out_trap_vector
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [31:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [31:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [31:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [31:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [31:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [31:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [31:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
  reg [31:0] _RAND_3350;
  reg [31:0] _RAND_3351;
  reg [31:0] _RAND_3352;
  reg [31:0] _RAND_3353;
  reg [31:0] _RAND_3354;
  reg [31:0] _RAND_3355;
  reg [31:0] _RAND_3356;
  reg [31:0] _RAND_3357;
  reg [31:0] _RAND_3358;
  reg [31:0] _RAND_3359;
  reg [31:0] _RAND_3360;
  reg [31:0] _RAND_3361;
  reg [31:0] _RAND_3362;
  reg [31:0] _RAND_3363;
  reg [31:0] _RAND_3364;
  reg [31:0] _RAND_3365;
  reg [31:0] _RAND_3366;
  reg [31:0] _RAND_3367;
  reg [31:0] _RAND_3368;
  reg [31:0] _RAND_3369;
  reg [31:0] _RAND_3370;
  reg [31:0] _RAND_3371;
  reg [31:0] _RAND_3372;
  reg [31:0] _RAND_3373;
  reg [31:0] _RAND_3374;
  reg [31:0] _RAND_3375;
  reg [31:0] _RAND_3376;
  reg [31:0] _RAND_3377;
  reg [31:0] _RAND_3378;
  reg [31:0] _RAND_3379;
  reg [31:0] _RAND_3380;
  reg [31:0] _RAND_3381;
  reg [31:0] _RAND_3382;
  reg [31:0] _RAND_3383;
  reg [31:0] _RAND_3384;
  reg [31:0] _RAND_3385;
  reg [31:0] _RAND_3386;
  reg [31:0] _RAND_3387;
  reg [31:0] _RAND_3388;
  reg [31:0] _RAND_3389;
  reg [31:0] _RAND_3390;
  reg [31:0] _RAND_3391;
  reg [31:0] _RAND_3392;
  reg [31:0] _RAND_3393;
  reg [31:0] _RAND_3394;
  reg [31:0] _RAND_3395;
  reg [31:0] _RAND_3396;
  reg [31:0] _RAND_3397;
  reg [31:0] _RAND_3398;
  reg [31:0] _RAND_3399;
  reg [31:0] _RAND_3400;
  reg [31:0] _RAND_3401;
  reg [31:0] _RAND_3402;
  reg [31:0] _RAND_3403;
  reg [31:0] _RAND_3404;
  reg [31:0] _RAND_3405;
  reg [31:0] _RAND_3406;
  reg [31:0] _RAND_3407;
  reg [31:0] _RAND_3408;
  reg [31:0] _RAND_3409;
  reg [31:0] _RAND_3410;
  reg [31:0] _RAND_3411;
  reg [31:0] _RAND_3412;
  reg [31:0] _RAND_3413;
  reg [31:0] _RAND_3414;
  reg [31:0] _RAND_3415;
  reg [31:0] _RAND_3416;
  reg [31:0] _RAND_3417;
  reg [31:0] _RAND_3418;
  reg [31:0] _RAND_3419;
  reg [31:0] _RAND_3420;
  reg [31:0] _RAND_3421;
  reg [31:0] _RAND_3422;
  reg [31:0] _RAND_3423;
  reg [31:0] _RAND_3424;
  reg [31:0] _RAND_3425;
  reg [31:0] _RAND_3426;
  reg [31:0] _RAND_3427;
  reg [31:0] _RAND_3428;
  reg [31:0] _RAND_3429;
  reg [31:0] _RAND_3430;
  reg [31:0] _RAND_3431;
  reg [31:0] _RAND_3432;
  reg [31:0] _RAND_3433;
  reg [31:0] _RAND_3434;
  reg [31:0] _RAND_3435;
  reg [31:0] _RAND_3436;
  reg [31:0] _RAND_3437;
  reg [31:0] _RAND_3438;
  reg [31:0] _RAND_3439;
  reg [31:0] _RAND_3440;
  reg [31:0] _RAND_3441;
  reg [31:0] _RAND_3442;
  reg [31:0] _RAND_3443;
  reg [31:0] _RAND_3444;
  reg [31:0] _RAND_3445;
  reg [31:0] _RAND_3446;
  reg [31:0] _RAND_3447;
  reg [31:0] _RAND_3448;
  reg [31:0] _RAND_3449;
  reg [31:0] _RAND_3450;
  reg [31:0] _RAND_3451;
  reg [31:0] _RAND_3452;
  reg [31:0] _RAND_3453;
  reg [31:0] _RAND_3454;
  reg [31:0] _RAND_3455;
  reg [31:0] _RAND_3456;
  reg [31:0] _RAND_3457;
  reg [31:0] _RAND_3458;
  reg [31:0] _RAND_3459;
  reg [31:0] _RAND_3460;
  reg [31:0] _RAND_3461;
  reg [31:0] _RAND_3462;
  reg [31:0] _RAND_3463;
  reg [31:0] _RAND_3464;
  reg [31:0] _RAND_3465;
  reg [31:0] _RAND_3466;
  reg [31:0] _RAND_3467;
  reg [31:0] _RAND_3468;
  reg [31:0] _RAND_3469;
  reg [31:0] _RAND_3470;
  reg [31:0] _RAND_3471;
  reg [31:0] _RAND_3472;
  reg [31:0] _RAND_3473;
  reg [31:0] _RAND_3474;
  reg [31:0] _RAND_3475;
  reg [31:0] _RAND_3476;
  reg [31:0] _RAND_3477;
  reg [31:0] _RAND_3478;
  reg [31:0] _RAND_3479;
  reg [31:0] _RAND_3480;
  reg [31:0] _RAND_3481;
  reg [31:0] _RAND_3482;
  reg [31:0] _RAND_3483;
  reg [31:0] _RAND_3484;
  reg [31:0] _RAND_3485;
  reg [31:0] _RAND_3486;
  reg [31:0] _RAND_3487;
  reg [31:0] _RAND_3488;
  reg [31:0] _RAND_3489;
  reg [31:0] _RAND_3490;
  reg [31:0] _RAND_3491;
  reg [31:0] _RAND_3492;
  reg [31:0] _RAND_3493;
  reg [31:0] _RAND_3494;
  reg [31:0] _RAND_3495;
  reg [31:0] _RAND_3496;
  reg [31:0] _RAND_3497;
  reg [31:0] _RAND_3498;
  reg [31:0] _RAND_3499;
  reg [31:0] _RAND_3500;
  reg [31:0] _RAND_3501;
  reg [31:0] _RAND_3502;
  reg [31:0] _RAND_3503;
  reg [31:0] _RAND_3504;
  reg [31:0] _RAND_3505;
  reg [31:0] _RAND_3506;
  reg [31:0] _RAND_3507;
  reg [31:0] _RAND_3508;
  reg [31:0] _RAND_3509;
  reg [31:0] _RAND_3510;
  reg [31:0] _RAND_3511;
  reg [31:0] _RAND_3512;
  reg [31:0] _RAND_3513;
  reg [31:0] _RAND_3514;
  reg [31:0] _RAND_3515;
  reg [31:0] _RAND_3516;
  reg [31:0] _RAND_3517;
  reg [31:0] _RAND_3518;
  reg [31:0] _RAND_3519;
  reg [31:0] _RAND_3520;
  reg [31:0] _RAND_3521;
  reg [31:0] _RAND_3522;
  reg [31:0] _RAND_3523;
  reg [31:0] _RAND_3524;
  reg [31:0] _RAND_3525;
  reg [31:0] _RAND_3526;
  reg [31:0] _RAND_3527;
  reg [31:0] _RAND_3528;
  reg [31:0] _RAND_3529;
  reg [31:0] _RAND_3530;
  reg [31:0] _RAND_3531;
  reg [31:0] _RAND_3532;
  reg [31:0] _RAND_3533;
  reg [31:0] _RAND_3534;
  reg [31:0] _RAND_3535;
  reg [31:0] _RAND_3536;
  reg [31:0] _RAND_3537;
  reg [31:0] _RAND_3538;
  reg [31:0] _RAND_3539;
  reg [31:0] _RAND_3540;
  reg [31:0] _RAND_3541;
  reg [31:0] _RAND_3542;
  reg [31:0] _RAND_3543;
  reg [31:0] _RAND_3544;
  reg [31:0] _RAND_3545;
  reg [31:0] _RAND_3546;
  reg [31:0] _RAND_3547;
  reg [31:0] _RAND_3548;
  reg [31:0] _RAND_3549;
  reg [31:0] _RAND_3550;
  reg [31:0] _RAND_3551;
  reg [31:0] _RAND_3552;
  reg [31:0] _RAND_3553;
  reg [31:0] _RAND_3554;
  reg [31:0] _RAND_3555;
  reg [31:0] _RAND_3556;
  reg [31:0] _RAND_3557;
  reg [31:0] _RAND_3558;
  reg [31:0] _RAND_3559;
  reg [31:0] _RAND_3560;
  reg [31:0] _RAND_3561;
  reg [31:0] _RAND_3562;
  reg [31:0] _RAND_3563;
  reg [31:0] _RAND_3564;
  reg [31:0] _RAND_3565;
  reg [31:0] _RAND_3566;
  reg [31:0] _RAND_3567;
  reg [31:0] _RAND_3568;
  reg [31:0] _RAND_3569;
  reg [31:0] _RAND_3570;
  reg [31:0] _RAND_3571;
  reg [31:0] _RAND_3572;
  reg [31:0] _RAND_3573;
  reg [31:0] _RAND_3574;
  reg [31:0] _RAND_3575;
  reg [31:0] _RAND_3576;
  reg [31:0] _RAND_3577;
  reg [31:0] _RAND_3578;
  reg [31:0] _RAND_3579;
  reg [31:0] _RAND_3580;
  reg [31:0] _RAND_3581;
  reg [31:0] _RAND_3582;
  reg [31:0] _RAND_3583;
  reg [31:0] _RAND_3584;
  reg [31:0] _RAND_3585;
  reg [31:0] _RAND_3586;
  reg [31:0] _RAND_3587;
  reg [31:0] _RAND_3588;
  reg [31:0] _RAND_3589;
  reg [31:0] _RAND_3590;
  reg [31:0] _RAND_3591;
  reg [31:0] _RAND_3592;
  reg [31:0] _RAND_3593;
  reg [31:0] _RAND_3594;
  reg [31:0] _RAND_3595;
  reg [31:0] _RAND_3596;
  reg [31:0] _RAND_3597;
  reg [31:0] _RAND_3598;
  reg [31:0] _RAND_3599;
  reg [31:0] _RAND_3600;
  reg [31:0] _RAND_3601;
  reg [31:0] _RAND_3602;
  reg [31:0] _RAND_3603;
  reg [31:0] _RAND_3604;
  reg [31:0] _RAND_3605;
  reg [31:0] _RAND_3606;
  reg [31:0] _RAND_3607;
  reg [31:0] _RAND_3608;
  reg [31:0] _RAND_3609;
  reg [31:0] _RAND_3610;
  reg [31:0] _RAND_3611;
  reg [31:0] _RAND_3612;
  reg [31:0] _RAND_3613;
  reg [31:0] _RAND_3614;
  reg [31:0] _RAND_3615;
  reg [31:0] _RAND_3616;
  reg [31:0] _RAND_3617;
  reg [31:0] _RAND_3618;
  reg [31:0] _RAND_3619;
  reg [31:0] _RAND_3620;
  reg [31:0] _RAND_3621;
  reg [31:0] _RAND_3622;
  reg [31:0] _RAND_3623;
  reg [31:0] _RAND_3624;
  reg [31:0] _RAND_3625;
  reg [31:0] _RAND_3626;
  reg [31:0] _RAND_3627;
  reg [31:0] _RAND_3628;
  reg [31:0] _RAND_3629;
  reg [31:0] _RAND_3630;
  reg [31:0] _RAND_3631;
  reg [31:0] _RAND_3632;
  reg [31:0] _RAND_3633;
  reg [31:0] _RAND_3634;
  reg [31:0] _RAND_3635;
  reg [31:0] _RAND_3636;
  reg [31:0] _RAND_3637;
  reg [31:0] _RAND_3638;
  reg [31:0] _RAND_3639;
  reg [31:0] _RAND_3640;
  reg [31:0] _RAND_3641;
  reg [31:0] _RAND_3642;
  reg [31:0] _RAND_3643;
  reg [31:0] _RAND_3644;
  reg [31:0] _RAND_3645;
  reg [31:0] _RAND_3646;
  reg [31:0] _RAND_3647;
  reg [31:0] _RAND_3648;
  reg [31:0] _RAND_3649;
  reg [31:0] _RAND_3650;
  reg [31:0] _RAND_3651;
  reg [31:0] _RAND_3652;
  reg [31:0] _RAND_3653;
  reg [31:0] _RAND_3654;
  reg [31:0] _RAND_3655;
  reg [31:0] _RAND_3656;
  reg [31:0] _RAND_3657;
  reg [31:0] _RAND_3658;
  reg [31:0] _RAND_3659;
  reg [31:0] _RAND_3660;
  reg [31:0] _RAND_3661;
  reg [31:0] _RAND_3662;
  reg [31:0] _RAND_3663;
  reg [31:0] _RAND_3664;
  reg [31:0] _RAND_3665;
  reg [31:0] _RAND_3666;
  reg [31:0] _RAND_3667;
  reg [31:0] _RAND_3668;
  reg [31:0] _RAND_3669;
  reg [31:0] _RAND_3670;
  reg [31:0] _RAND_3671;
  reg [31:0] _RAND_3672;
  reg [31:0] _RAND_3673;
  reg [31:0] _RAND_3674;
  reg [31:0] _RAND_3675;
  reg [31:0] _RAND_3676;
  reg [31:0] _RAND_3677;
  reg [31:0] _RAND_3678;
  reg [31:0] _RAND_3679;
  reg [31:0] _RAND_3680;
  reg [31:0] _RAND_3681;
  reg [31:0] _RAND_3682;
  reg [31:0] _RAND_3683;
  reg [31:0] _RAND_3684;
  reg [31:0] _RAND_3685;
  reg [31:0] _RAND_3686;
  reg [31:0] _RAND_3687;
  reg [31:0] _RAND_3688;
  reg [31:0] _RAND_3689;
  reg [31:0] _RAND_3690;
  reg [31:0] _RAND_3691;
  reg [31:0] _RAND_3692;
  reg [31:0] _RAND_3693;
  reg [31:0] _RAND_3694;
  reg [31:0] _RAND_3695;
  reg [31:0] _RAND_3696;
  reg [31:0] _RAND_3697;
  reg [31:0] _RAND_3698;
  reg [31:0] _RAND_3699;
  reg [31:0] _RAND_3700;
  reg [31:0] _RAND_3701;
  reg [31:0] _RAND_3702;
  reg [31:0] _RAND_3703;
  reg [31:0] _RAND_3704;
  reg [31:0] _RAND_3705;
  reg [31:0] _RAND_3706;
  reg [31:0] _RAND_3707;
  reg [31:0] _RAND_3708;
  reg [31:0] _RAND_3709;
  reg [31:0] _RAND_3710;
  reg [31:0] _RAND_3711;
  reg [31:0] _RAND_3712;
  reg [31:0] _RAND_3713;
  reg [31:0] _RAND_3714;
  reg [31:0] _RAND_3715;
  reg [31:0] _RAND_3716;
  reg [31:0] _RAND_3717;
  reg [31:0] _RAND_3718;
  reg [31:0] _RAND_3719;
  reg [31:0] _RAND_3720;
  reg [31:0] _RAND_3721;
  reg [31:0] _RAND_3722;
  reg [31:0] _RAND_3723;
  reg [31:0] _RAND_3724;
  reg [31:0] _RAND_3725;
  reg [31:0] _RAND_3726;
  reg [31:0] _RAND_3727;
  reg [31:0] _RAND_3728;
  reg [31:0] _RAND_3729;
  reg [31:0] _RAND_3730;
  reg [31:0] _RAND_3731;
  reg [31:0] _RAND_3732;
  reg [31:0] _RAND_3733;
  reg [31:0] _RAND_3734;
  reg [31:0] _RAND_3735;
  reg [31:0] _RAND_3736;
  reg [31:0] _RAND_3737;
  reg [31:0] _RAND_3738;
  reg [31:0] _RAND_3739;
  reg [31:0] _RAND_3740;
  reg [31:0] _RAND_3741;
  reg [31:0] _RAND_3742;
  reg [31:0] _RAND_3743;
  reg [31:0] _RAND_3744;
  reg [31:0] _RAND_3745;
  reg [31:0] _RAND_3746;
  reg [31:0] _RAND_3747;
  reg [31:0] _RAND_3748;
  reg [31:0] _RAND_3749;
  reg [31:0] _RAND_3750;
  reg [31:0] _RAND_3751;
  reg [31:0] _RAND_3752;
  reg [31:0] _RAND_3753;
  reg [31:0] _RAND_3754;
  reg [31:0] _RAND_3755;
  reg [31:0] _RAND_3756;
  reg [31:0] _RAND_3757;
  reg [31:0] _RAND_3758;
  reg [31:0] _RAND_3759;
  reg [31:0] _RAND_3760;
  reg [31:0] _RAND_3761;
  reg [31:0] _RAND_3762;
  reg [31:0] _RAND_3763;
  reg [31:0] _RAND_3764;
  reg [31:0] _RAND_3765;
  reg [31:0] _RAND_3766;
  reg [31:0] _RAND_3767;
  reg [31:0] _RAND_3768;
  reg [31:0] _RAND_3769;
  reg [31:0] _RAND_3770;
  reg [31:0] _RAND_3771;
  reg [31:0] _RAND_3772;
  reg [31:0] _RAND_3773;
  reg [31:0] _RAND_3774;
  reg [31:0] _RAND_3775;
  reg [31:0] _RAND_3776;
  reg [31:0] _RAND_3777;
  reg [31:0] _RAND_3778;
  reg [31:0] _RAND_3779;
  reg [31:0] _RAND_3780;
  reg [31:0] _RAND_3781;
  reg [31:0] _RAND_3782;
  reg [31:0] _RAND_3783;
  reg [31:0] _RAND_3784;
  reg [31:0] _RAND_3785;
  reg [31:0] _RAND_3786;
  reg [31:0] _RAND_3787;
  reg [31:0] _RAND_3788;
  reg [31:0] _RAND_3789;
  reg [31:0] _RAND_3790;
  reg [31:0] _RAND_3791;
  reg [31:0] _RAND_3792;
  reg [31:0] _RAND_3793;
  reg [31:0] _RAND_3794;
  reg [31:0] _RAND_3795;
  reg [31:0] _RAND_3796;
  reg [31:0] _RAND_3797;
  reg [31:0] _RAND_3798;
  reg [31:0] _RAND_3799;
  reg [31:0] _RAND_3800;
  reg [31:0] _RAND_3801;
  reg [31:0] _RAND_3802;
  reg [31:0] _RAND_3803;
  reg [31:0] _RAND_3804;
  reg [31:0] _RAND_3805;
  reg [31:0] _RAND_3806;
  reg [31:0] _RAND_3807;
  reg [31:0] _RAND_3808;
  reg [31:0] _RAND_3809;
  reg [31:0] _RAND_3810;
  reg [31:0] _RAND_3811;
  reg [31:0] _RAND_3812;
  reg [31:0] _RAND_3813;
  reg [31:0] _RAND_3814;
  reg [31:0] _RAND_3815;
  reg [31:0] _RAND_3816;
  reg [31:0] _RAND_3817;
  reg [31:0] _RAND_3818;
  reg [31:0] _RAND_3819;
  reg [31:0] _RAND_3820;
  reg [31:0] _RAND_3821;
  reg [31:0] _RAND_3822;
  reg [31:0] _RAND_3823;
  reg [31:0] _RAND_3824;
  reg [31:0] _RAND_3825;
  reg [31:0] _RAND_3826;
  reg [31:0] _RAND_3827;
  reg [31:0] _RAND_3828;
  reg [31:0] _RAND_3829;
  reg [31:0] _RAND_3830;
  reg [31:0] _RAND_3831;
  reg [31:0] _RAND_3832;
  reg [31:0] _RAND_3833;
  reg [31:0] _RAND_3834;
  reg [31:0] _RAND_3835;
  reg [31:0] _RAND_3836;
  reg [31:0] _RAND_3837;
  reg [31:0] _RAND_3838;
  reg [31:0] _RAND_3839;
  reg [31:0] _RAND_3840;
  reg [31:0] _RAND_3841;
  reg [31:0] _RAND_3842;
  reg [31:0] _RAND_3843;
  reg [31:0] _RAND_3844;
  reg [31:0] _RAND_3845;
  reg [31:0] _RAND_3846;
  reg [31:0] _RAND_3847;
  reg [31:0] _RAND_3848;
  reg [31:0] _RAND_3849;
  reg [31:0] _RAND_3850;
  reg [31:0] _RAND_3851;
  reg [31:0] _RAND_3852;
  reg [31:0] _RAND_3853;
  reg [31:0] _RAND_3854;
  reg [31:0] _RAND_3855;
  reg [31:0] _RAND_3856;
  reg [31:0] _RAND_3857;
  reg [31:0] _RAND_3858;
  reg [31:0] _RAND_3859;
  reg [31:0] _RAND_3860;
  reg [31:0] _RAND_3861;
  reg [31:0] _RAND_3862;
  reg [31:0] _RAND_3863;
  reg [31:0] _RAND_3864;
  reg [31:0] _RAND_3865;
  reg [31:0] _RAND_3866;
  reg [31:0] _RAND_3867;
  reg [31:0] _RAND_3868;
  reg [31:0] _RAND_3869;
  reg [31:0] _RAND_3870;
  reg [31:0] _RAND_3871;
  reg [31:0] _RAND_3872;
  reg [31:0] _RAND_3873;
  reg [31:0] _RAND_3874;
  reg [31:0] _RAND_3875;
  reg [31:0] _RAND_3876;
  reg [31:0] _RAND_3877;
  reg [31:0] _RAND_3878;
  reg [31:0] _RAND_3879;
  reg [31:0] _RAND_3880;
  reg [31:0] _RAND_3881;
  reg [31:0] _RAND_3882;
  reg [31:0] _RAND_3883;
  reg [31:0] _RAND_3884;
  reg [31:0] _RAND_3885;
  reg [31:0] _RAND_3886;
  reg [31:0] _RAND_3887;
  reg [31:0] _RAND_3888;
  reg [31:0] _RAND_3889;
  reg [31:0] _RAND_3890;
  reg [31:0] _RAND_3891;
  reg [31:0] _RAND_3892;
  reg [31:0] _RAND_3893;
  reg [31:0] _RAND_3894;
  reg [31:0] _RAND_3895;
  reg [31:0] _RAND_3896;
  reg [31:0] _RAND_3897;
  reg [31:0] _RAND_3898;
  reg [31:0] _RAND_3899;
  reg [31:0] _RAND_3900;
  reg [31:0] _RAND_3901;
  reg [31:0] _RAND_3902;
  reg [31:0] _RAND_3903;
  reg [31:0] _RAND_3904;
  reg [31:0] _RAND_3905;
  reg [31:0] _RAND_3906;
  reg [31:0] _RAND_3907;
  reg [31:0] _RAND_3908;
  reg [31:0] _RAND_3909;
  reg [31:0] _RAND_3910;
  reg [31:0] _RAND_3911;
  reg [31:0] _RAND_3912;
  reg [31:0] _RAND_3913;
  reg [31:0] _RAND_3914;
  reg [31:0] _RAND_3915;
  reg [31:0] _RAND_3916;
  reg [31:0] _RAND_3917;
  reg [31:0] _RAND_3918;
  reg [31:0] _RAND_3919;
  reg [31:0] _RAND_3920;
  reg [31:0] _RAND_3921;
  reg [31:0] _RAND_3922;
  reg [31:0] _RAND_3923;
  reg [31:0] _RAND_3924;
  reg [31:0] _RAND_3925;
  reg [31:0] _RAND_3926;
  reg [31:0] _RAND_3927;
  reg [31:0] _RAND_3928;
  reg [31:0] _RAND_3929;
  reg [31:0] _RAND_3930;
  reg [31:0] _RAND_3931;
  reg [31:0] _RAND_3932;
  reg [31:0] _RAND_3933;
  reg [31:0] _RAND_3934;
  reg [31:0] _RAND_3935;
  reg [31:0] _RAND_3936;
  reg [31:0] _RAND_3937;
  reg [31:0] _RAND_3938;
  reg [31:0] _RAND_3939;
  reg [31:0] _RAND_3940;
  reg [31:0] _RAND_3941;
  reg [31:0] _RAND_3942;
  reg [31:0] _RAND_3943;
  reg [31:0] _RAND_3944;
  reg [31:0] _RAND_3945;
  reg [31:0] _RAND_3946;
  reg [31:0] _RAND_3947;
  reg [31:0] _RAND_3948;
  reg [31:0] _RAND_3949;
  reg [31:0] _RAND_3950;
  reg [31:0] _RAND_3951;
  reg [31:0] _RAND_3952;
  reg [31:0] _RAND_3953;
  reg [31:0] _RAND_3954;
  reg [31:0] _RAND_3955;
  reg [31:0] _RAND_3956;
  reg [31:0] _RAND_3957;
  reg [31:0] _RAND_3958;
  reg [31:0] _RAND_3959;
  reg [31:0] _RAND_3960;
  reg [31:0] _RAND_3961;
  reg [31:0] _RAND_3962;
  reg [31:0] _RAND_3963;
  reg [31:0] _RAND_3964;
  reg [31:0] _RAND_3965;
  reg [31:0] _RAND_3966;
  reg [31:0] _RAND_3967;
  reg [31:0] _RAND_3968;
  reg [31:0] _RAND_3969;
  reg [31:0] _RAND_3970;
  reg [31:0] _RAND_3971;
  reg [31:0] _RAND_3972;
  reg [31:0] _RAND_3973;
  reg [31:0] _RAND_3974;
  reg [31:0] _RAND_3975;
  reg [31:0] _RAND_3976;
  reg [31:0] _RAND_3977;
  reg [31:0] _RAND_3978;
  reg [31:0] _RAND_3979;
  reg [31:0] _RAND_3980;
  reg [31:0] _RAND_3981;
  reg [31:0] _RAND_3982;
  reg [31:0] _RAND_3983;
  reg [31:0] _RAND_3984;
  reg [31:0] _RAND_3985;
  reg [31:0] _RAND_3986;
  reg [31:0] _RAND_3987;
  reg [31:0] _RAND_3988;
  reg [31:0] _RAND_3989;
  reg [31:0] _RAND_3990;
  reg [31:0] _RAND_3991;
  reg [31:0] _RAND_3992;
  reg [31:0] _RAND_3993;
  reg [31:0] _RAND_3994;
  reg [31:0] _RAND_3995;
  reg [31:0] _RAND_3996;
  reg [31:0] _RAND_3997;
  reg [31:0] _RAND_3998;
  reg [31:0] _RAND_3999;
  reg [31:0] _RAND_4000;
  reg [31:0] _RAND_4001;
  reg [31:0] _RAND_4002;
  reg [31:0] _RAND_4003;
  reg [31:0] _RAND_4004;
  reg [31:0] _RAND_4005;
  reg [31:0] _RAND_4006;
  reg [31:0] _RAND_4007;
  reg [31:0] _RAND_4008;
  reg [31:0] _RAND_4009;
  reg [31:0] _RAND_4010;
  reg [31:0] _RAND_4011;
  reg [31:0] _RAND_4012;
  reg [31:0] _RAND_4013;
  reg [31:0] _RAND_4014;
  reg [31:0] _RAND_4015;
  reg [31:0] _RAND_4016;
  reg [31:0] _RAND_4017;
  reg [31:0] _RAND_4018;
  reg [31:0] _RAND_4019;
  reg [31:0] _RAND_4020;
  reg [31:0] _RAND_4021;
  reg [31:0] _RAND_4022;
  reg [31:0] _RAND_4023;
  reg [31:0] _RAND_4024;
  reg [31:0] _RAND_4025;
  reg [31:0] _RAND_4026;
  reg [31:0] _RAND_4027;
  reg [31:0] _RAND_4028;
  reg [31:0] _RAND_4029;
  reg [31:0] _RAND_4030;
  reg [31:0] _RAND_4031;
  reg [31:0] _RAND_4032;
  reg [31:0] _RAND_4033;
  reg [31:0] _RAND_4034;
  reg [31:0] _RAND_4035;
  reg [31:0] _RAND_4036;
  reg [31:0] _RAND_4037;
  reg [31:0] _RAND_4038;
  reg [31:0] _RAND_4039;
  reg [31:0] _RAND_4040;
  reg [31:0] _RAND_4041;
  reg [31:0] _RAND_4042;
  reg [31:0] _RAND_4043;
  reg [31:0] _RAND_4044;
  reg [31:0] _RAND_4045;
  reg [31:0] _RAND_4046;
  reg [31:0] _RAND_4047;
  reg [31:0] _RAND_4048;
  reg [31:0] _RAND_4049;
  reg [31:0] _RAND_4050;
  reg [31:0] _RAND_4051;
  reg [31:0] _RAND_4052;
  reg [31:0] _RAND_4053;
  reg [31:0] _RAND_4054;
  reg [31:0] _RAND_4055;
  reg [31:0] _RAND_4056;
  reg [31:0] _RAND_4057;
  reg [31:0] _RAND_4058;
  reg [31:0] _RAND_4059;
  reg [31:0] _RAND_4060;
  reg [31:0] _RAND_4061;
  reg [31:0] _RAND_4062;
  reg [31:0] _RAND_4063;
  reg [31:0] _RAND_4064;
  reg [31:0] _RAND_4065;
  reg [31:0] _RAND_4066;
  reg [31:0] _RAND_4067;
  reg [31:0] _RAND_4068;
  reg [31:0] _RAND_4069;
  reg [31:0] _RAND_4070;
  reg [31:0] _RAND_4071;
  reg [31:0] _RAND_4072;
  reg [31:0] _RAND_4073;
  reg [31:0] _RAND_4074;
  reg [31:0] _RAND_4075;
  reg [31:0] _RAND_4076;
  reg [31:0] _RAND_4077;
  reg [31:0] _RAND_4078;
  reg [31:0] _RAND_4079;
  reg [31:0] _RAND_4080;
  reg [31:0] _RAND_4081;
  reg [31:0] _RAND_4082;
  reg [31:0] _RAND_4083;
  reg [31:0] _RAND_4084;
  reg [31:0] _RAND_4085;
  reg [31:0] _RAND_4086;
  reg [31:0] _RAND_4087;
  reg [31:0] _RAND_4088;
  reg [31:0] _RAND_4089;
  reg [31:0] _RAND_4090;
  reg [31:0] _RAND_4091;
  reg [31:0] _RAND_4092;
  reg [31:0] _RAND_4093;
  reg [31:0] _RAND_4094;
  reg [31:0] _RAND_4095;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_csr_0; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_5; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_6; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_7; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_8; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_9; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_10; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_11; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_12; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_13; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_14; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_15; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_16; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_17; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_18; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_19; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_20; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_21; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_22; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_23; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_24; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_25; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_26; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_27; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_28; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_29; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_30; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_31; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_32; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_33; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_34; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_35; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_36; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_37; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_38; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_39; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_40; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_41; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_42; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_43; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_44; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_45; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_46; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_47; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_48; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_49; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_50; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_51; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_52; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_53; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_54; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_55; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_56; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_57; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_58; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_59; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_60; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_61; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_62; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_63; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_64; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_65; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_66; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_67; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_68; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_69; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_70; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_71; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_72; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_73; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_74; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_75; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_76; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_77; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_78; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_79; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_80; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_81; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_82; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_83; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_84; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_85; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_86; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_87; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_88; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_89; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_90; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_91; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_92; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_93; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_94; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_95; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_96; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_97; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_98; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_99; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_100; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_101; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_102; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_103; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_104; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_105; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_106; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_107; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_108; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_109; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_110; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_111; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_112; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_113; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_114; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_115; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_116; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_117; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_118; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_119; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_120; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_121; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_122; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_123; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_124; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_125; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_126; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_127; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_128; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_129; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_130; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_131; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_132; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_133; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_134; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_135; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_136; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_137; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_138; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_139; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_140; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_141; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_142; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_143; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_144; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_145; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_146; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_147; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_148; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_149; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_150; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_151; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_152; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_153; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_154; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_155; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_156; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_157; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_158; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_159; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_160; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_161; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_162; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_163; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_164; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_165; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_166; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_167; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_168; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_169; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_170; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_171; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_172; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_173; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_174; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_175; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_176; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_177; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_178; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_179; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_180; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_181; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_182; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_183; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_184; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_185; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_186; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_187; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_188; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_189; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_190; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_191; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_192; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_193; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_194; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_195; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_196; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_197; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_198; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_199; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_200; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_201; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_202; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_203; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_204; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_205; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_206; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_207; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_208; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_209; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_210; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_211; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_212; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_213; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_214; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_215; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_216; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_217; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_218; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_219; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_220; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_221; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_222; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_223; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_224; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_225; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_226; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_227; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_228; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_229; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_230; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_231; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_232; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_233; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_234; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_235; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_236; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_237; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_238; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_239; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_240; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_241; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_242; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_243; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_244; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_245; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_246; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_247; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_248; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_249; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_250; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_251; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_252; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_253; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_254; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_255; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_256; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_257; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_258; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_259; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_260; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_261; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_262; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_263; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_264; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_265; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_266; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_267; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_268; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_269; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_270; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_271; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_272; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_273; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_274; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_275; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_276; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_277; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_278; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_279; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_280; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_281; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_282; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_283; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_284; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_285; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_286; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_287; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_288; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_289; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_290; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_291; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_292; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_293; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_294; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_295; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_296; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_297; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_298; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_299; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_300; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_301; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_302; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_303; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_304; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_305; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_306; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_307; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_308; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_309; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_310; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_311; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_312; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_313; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_314; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_315; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_316; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_317; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_318; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_319; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_320; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_321; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_322; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_323; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_324; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_325; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_326; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_327; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_328; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_329; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_330; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_331; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_332; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_333; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_334; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_335; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_336; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_337; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_338; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_339; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_340; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_341; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_342; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_343; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_344; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_345; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_346; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_347; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_348; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_349; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_350; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_351; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_352; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_353; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_354; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_355; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_356; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_357; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_358; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_359; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_360; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_361; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_362; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_363; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_364; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_365; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_366; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_367; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_368; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_369; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_370; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_371; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_372; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_373; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_374; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_375; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_376; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_377; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_378; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_379; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_380; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_381; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_382; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_383; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_384; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_385; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_386; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_387; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_388; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_389; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_390; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_391; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_392; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_393; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_394; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_395; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_396; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_397; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_398; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_399; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_400; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_401; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_402; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_403; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_404; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_405; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_406; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_407; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_408; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_409; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_410; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_411; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_412; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_413; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_414; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_415; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_416; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_417; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_418; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_419; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_420; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_421; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_422; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_423; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_424; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_425; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_426; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_427; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_428; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_429; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_430; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_431; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_432; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_433; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_434; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_435; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_436; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_437; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_438; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_439; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_440; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_441; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_442; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_443; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_444; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_445; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_446; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_447; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_448; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_449; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_450; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_451; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_452; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_453; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_454; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_455; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_456; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_457; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_458; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_459; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_460; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_461; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_462; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_463; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_464; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_465; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_466; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_467; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_468; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_469; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_470; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_471; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_472; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_473; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_474; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_475; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_476; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_477; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_478; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_479; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_480; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_481; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_482; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_483; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_484; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_485; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_486; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_487; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_488; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_489; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_490; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_491; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_492; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_493; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_494; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_495; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_496; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_497; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_498; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_499; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_500; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_501; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_502; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_503; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_504; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_505; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_506; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_507; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_508; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_509; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_510; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_511; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_512; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_513; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_514; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_515; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_516; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_517; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_518; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_519; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_520; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_521; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_522; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_523; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_524; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_525; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_526; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_527; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_528; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_529; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_530; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_531; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_532; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_533; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_534; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_535; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_536; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_537; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_538; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_539; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_540; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_541; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_542; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_543; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_544; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_545; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_546; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_547; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_548; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_549; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_550; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_551; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_552; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_553; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_554; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_555; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_556; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_557; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_558; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_559; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_560; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_561; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_562; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_563; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_564; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_565; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_566; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_567; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_568; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_569; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_570; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_571; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_572; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_573; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_574; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_575; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_576; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_577; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_578; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_579; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_580; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_581; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_582; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_583; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_584; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_585; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_586; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_587; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_588; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_589; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_590; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_591; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_592; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_593; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_594; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_595; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_596; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_597; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_598; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_599; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_600; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_601; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_602; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_603; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_604; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_605; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_606; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_607; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_608; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_609; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_610; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_611; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_612; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_613; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_614; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_615; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_616; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_617; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_618; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_619; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_620; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_621; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_622; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_623; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_624; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_625; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_626; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_627; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_628; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_629; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_630; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_631; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_632; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_633; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_634; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_635; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_636; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_637; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_638; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_639; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_640; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_641; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_642; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_643; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_644; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_645; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_646; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_647; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_648; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_649; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_650; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_651; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_652; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_653; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_654; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_655; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_656; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_657; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_658; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_659; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_660; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_661; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_662; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_663; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_664; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_665; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_666; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_667; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_668; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_669; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_670; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_671; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_672; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_673; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_674; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_675; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_676; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_677; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_678; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_679; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_680; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_681; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_682; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_683; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_684; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_685; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_686; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_687; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_688; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_689; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_690; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_691; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_692; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_693; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_694; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_695; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_696; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_697; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_698; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_699; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_700; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_701; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_702; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_703; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_704; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_705; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_706; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_707; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_708; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_709; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_710; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_711; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_712; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_713; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_714; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_715; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_716; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_717; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_718; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_719; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_720; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_721; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_722; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_723; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_724; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_725; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_726; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_727; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_728; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_729; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_730; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_731; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_732; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_733; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_734; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_735; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_736; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_737; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_738; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_739; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_740; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_741; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_742; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_743; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_744; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_745; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_746; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_747; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_748; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_749; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_750; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_751; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_752; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_753; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_754; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_755; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_756; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_757; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_758; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_759; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_760; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_761; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_762; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_763; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_764; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_765; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_766; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_767; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_768; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_769; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_770; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_771; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_772; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_773; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_774; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_775; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_776; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_777; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_778; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_779; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_780; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_781; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_782; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_783; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_784; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_785; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_786; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_787; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_788; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_789; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_790; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_791; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_792; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_793; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_794; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_795; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_796; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_797; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_798; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_799; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_800; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_801; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_802; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_803; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_804; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_805; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_806; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_807; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_808; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_809; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_810; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_811; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_812; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_813; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_814; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_815; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_816; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_817; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_818; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_819; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_820; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_821; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_822; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_823; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_824; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_825; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_826; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_827; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_828; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_829; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_830; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_831; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_832; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_833; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_834; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_835; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_836; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_837; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_838; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_839; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_840; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_841; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_842; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_843; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_844; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_845; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_846; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_847; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_848; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_849; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_850; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_851; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_852; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_853; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_854; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_855; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_856; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_857; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_858; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_859; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_860; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_861; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_862; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_863; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_864; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_865; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_866; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_867; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_868; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_869; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_870; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_871; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_872; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_873; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_874; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_875; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_876; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_877; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_878; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_879; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_880; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_881; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_882; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_883; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_884; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_885; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_886; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_887; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_888; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_889; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_890; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_891; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_892; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_893; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_894; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_895; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_896; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_897; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_898; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_899; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_900; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_901; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_902; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_903; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_904; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_905; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_906; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_907; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_908; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_909; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_910; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_911; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_912; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_913; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_914; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_915; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_916; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_917; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_918; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_919; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_920; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_921; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_922; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_923; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_924; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_925; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_926; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_927; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_928; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_929; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_930; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_931; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_932; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_933; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_934; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_935; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_936; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_937; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_938; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_939; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_940; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_941; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_942; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_943; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_944; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_945; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_946; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_947; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_948; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_949; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_950; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_951; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_952; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_953; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_954; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_955; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_956; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_957; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_958; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_959; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_960; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_961; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_962; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_963; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_964; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_965; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_966; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_967; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_968; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_969; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_970; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_971; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_972; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_973; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_974; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_975; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_976; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_977; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_978; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_979; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_980; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_981; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_982; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_983; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_984; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_985; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_986; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_987; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_988; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_989; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_990; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_991; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_992; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_993; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_994; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_995; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_996; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_997; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_998; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_999; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1000; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1001; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1002; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1003; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1004; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1005; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1006; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1007; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1008; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1009; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1010; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1011; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1012; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1013; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1014; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1015; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1016; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1017; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1018; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1019; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1020; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1021; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1022; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1023; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1024; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1025; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1026; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1027; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1028; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1029; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1030; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1031; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1032; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1033; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1034; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1035; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1036; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1037; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1038; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1039; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1040; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1041; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1042; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1043; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1044; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1045; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1046; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1047; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1048; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1049; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1050; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1051; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1052; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1053; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1054; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1055; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1056; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1057; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1058; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1059; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1060; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1061; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1062; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1063; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1064; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1065; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1066; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1067; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1068; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1069; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1070; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1071; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1072; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1073; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1074; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1075; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1076; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1077; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1078; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1079; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1080; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1081; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1082; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1083; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1084; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1085; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1086; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1087; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1088; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1089; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1090; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1091; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1092; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1093; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1094; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1095; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1096; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1097; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1098; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1099; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1100; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1101; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1102; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1103; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1104; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1105; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1106; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1107; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1108; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1109; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1110; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1111; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1112; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1113; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1114; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1115; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1116; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1117; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1118; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1119; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1120; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1121; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1122; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1123; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1124; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1125; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1126; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1127; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1128; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1129; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1130; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1131; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1132; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1133; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1134; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1135; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1136; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1137; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1138; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1139; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1140; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1141; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1142; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1143; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1144; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1145; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1146; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1147; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1148; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1149; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1150; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1151; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1152; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1153; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1154; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1155; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1156; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1157; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1158; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1159; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1160; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1161; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1162; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1163; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1164; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1165; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1166; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1167; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1168; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1169; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1170; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1171; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1172; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1173; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1174; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1175; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1176; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1177; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1178; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1179; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1180; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1181; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1182; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1183; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1184; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1185; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1186; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1187; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1188; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1189; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1190; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1191; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1192; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1193; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1194; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1195; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1196; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1197; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1198; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1199; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1200; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1201; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1202; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1203; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1204; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1205; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1206; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1207; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1208; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1209; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1210; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1211; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1212; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1213; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1214; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1215; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1216; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1217; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1218; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1219; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1220; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1221; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1222; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1223; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1224; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1225; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1226; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1227; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1228; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1229; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1230; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1231; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1232; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1233; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1234; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1235; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1236; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1237; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1238; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1239; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1240; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1241; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1242; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1243; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1244; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1245; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1246; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1247; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1248; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1249; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1250; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1251; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1252; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1253; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1254; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1255; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1256; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1257; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1258; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1259; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1260; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1261; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1262; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1263; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1264; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1265; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1266; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1267; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1268; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1269; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1270; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1271; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1272; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1273; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1274; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1275; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1276; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1277; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1278; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1279; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1280; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1281; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1282; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1283; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1284; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1285; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1286; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1287; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1288; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1289; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1290; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1291; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1292; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1293; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1294; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1295; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1296; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1297; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1298; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1299; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1300; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1301; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1302; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1303; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1304; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1305; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1306; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1307; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1308; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1309; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1310; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1311; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1312; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1313; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1314; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1315; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1316; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1317; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1318; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1319; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1320; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1321; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1322; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1323; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1324; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1325; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1326; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1327; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1328; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1329; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1330; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1331; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1332; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1333; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1334; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1335; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1336; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1337; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1338; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1339; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1340; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1341; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1342; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1343; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1344; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1345; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1346; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1347; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1348; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1349; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1350; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1351; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1352; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1353; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1354; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1355; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1356; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1357; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1358; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1359; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1360; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1361; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1362; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1363; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1364; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1365; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1366; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1367; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1368; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1369; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1370; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1371; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1372; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1373; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1374; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1375; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1376; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1377; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1378; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1379; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1380; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1381; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1382; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1383; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1384; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1385; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1386; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1387; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1388; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1389; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1390; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1391; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1392; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1393; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1394; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1395; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1396; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1397; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1398; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1399; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1400; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1401; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1402; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1403; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1404; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1405; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1406; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1407; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1408; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1409; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1410; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1411; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1412; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1413; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1414; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1415; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1416; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1417; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1418; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1419; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1420; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1421; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1422; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1423; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1424; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1425; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1426; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1427; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1428; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1429; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1430; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1431; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1432; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1433; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1434; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1435; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1436; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1437; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1438; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1439; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1440; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1441; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1442; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1443; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1444; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1445; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1446; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1447; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1448; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1449; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1450; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1451; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1452; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1453; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1454; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1455; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1456; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1457; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1458; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1459; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1460; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1461; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1462; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1463; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1464; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1465; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1466; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1467; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1468; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1469; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1470; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1471; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1472; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1473; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1474; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1475; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1476; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1477; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1478; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1479; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1480; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1481; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1482; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1483; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1484; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1485; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1486; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1487; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1488; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1489; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1490; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1491; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1492; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1493; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1494; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1495; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1496; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1497; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1498; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1499; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1500; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1501; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1502; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1503; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1504; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1505; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1506; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1507; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1508; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1509; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1510; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1511; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1512; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1513; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1514; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1515; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1516; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1517; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1518; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1519; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1520; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1521; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1522; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1523; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1524; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1525; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1526; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1527; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1528; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1529; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1530; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1531; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1532; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1533; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1534; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1535; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1536; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1537; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1538; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1539; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1540; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1541; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1542; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1543; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1544; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1545; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1546; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1547; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1548; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1549; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1550; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1551; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1552; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1553; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1554; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1555; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1556; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1557; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1558; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1559; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1560; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1561; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1562; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1563; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1564; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1565; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1566; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1567; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1568; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1569; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1570; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1571; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1572; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1573; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1574; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1575; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1576; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1577; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1578; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1579; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1580; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1581; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1582; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1583; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1584; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1585; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1586; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1587; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1588; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1589; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1590; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1591; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1592; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1593; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1594; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1595; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1596; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1597; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1598; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1599; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1600; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1601; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1602; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1603; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1604; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1605; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1606; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1607; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1608; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1609; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1610; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1611; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1612; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1613; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1614; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1615; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1616; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1617; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1618; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1619; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1620; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1621; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1622; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1623; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1624; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1625; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1626; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1627; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1628; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1629; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1630; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1631; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1632; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1633; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1634; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1635; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1636; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1637; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1638; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1639; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1640; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1641; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1642; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1643; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1644; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1645; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1646; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1647; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1648; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1649; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1650; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1651; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1652; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1653; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1654; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1655; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1656; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1657; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1658; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1659; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1660; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1661; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1662; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1663; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1664; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1665; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1666; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1667; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1668; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1669; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1670; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1671; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1672; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1673; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1674; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1675; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1676; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1677; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1678; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1679; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1680; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1681; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1682; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1683; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1684; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1685; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1686; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1687; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1688; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1689; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1690; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1691; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1692; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1693; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1694; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1695; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1696; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1697; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1698; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1699; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1700; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1701; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1702; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1703; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1704; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1705; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1706; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1707; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1708; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1709; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1710; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1711; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1712; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1713; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1714; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1715; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1716; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1717; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1718; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1719; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1720; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1721; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1722; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1723; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1724; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1725; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1726; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1727; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1728; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1729; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1730; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1731; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1732; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1733; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1734; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1735; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1736; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1737; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1738; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1739; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1740; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1741; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1742; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1743; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1744; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1745; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1746; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1747; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1748; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1749; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1750; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1751; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1752; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1753; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1754; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1755; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1756; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1757; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1758; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1759; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1760; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1761; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1762; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1763; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1764; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1765; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1766; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1767; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1768; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1769; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1770; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1771; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1772; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1773; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1774; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1775; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1776; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1777; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1778; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1779; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1780; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1781; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1782; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1783; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1784; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1785; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1786; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1787; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1788; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1789; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1790; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1791; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1792; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1793; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1794; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1795; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1796; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1797; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1798; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1799; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1800; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1801; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1802; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1803; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1804; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1805; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1806; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1807; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1808; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1809; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1810; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1811; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1812; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1813; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1814; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1815; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1816; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1817; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1818; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1819; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1820; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1821; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1822; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1823; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1824; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1825; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1826; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1827; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1828; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1829; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1830; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1831; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1832; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1833; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1834; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1835; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1836; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1837; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1838; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1839; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1840; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1841; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1842; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1843; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1844; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1845; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1846; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1847; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1848; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1849; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1850; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1851; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1852; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1853; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1854; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1855; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1856; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1857; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1858; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1859; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1860; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1861; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1862; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1863; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1864; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1865; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1866; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1867; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1868; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1869; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1870; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1871; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1872; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1873; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1874; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1875; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1876; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1877; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1878; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1879; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1880; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1881; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1882; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1883; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1884; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1885; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1886; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1887; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1888; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1889; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1890; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1891; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1892; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1893; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1894; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1895; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1896; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1897; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1898; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1899; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1900; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1901; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1902; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1903; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1904; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1905; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1906; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1907; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1908; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1909; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1910; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1911; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1912; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1913; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1914; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1915; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1916; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1917; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1918; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1919; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1920; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1921; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1922; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1923; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1924; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1925; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1926; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1927; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1928; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1929; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1930; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1931; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1932; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1933; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1934; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1935; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1936; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1937; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1938; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1939; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1940; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1941; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1942; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1943; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1944; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1945; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1946; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1947; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1948; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1949; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1950; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1951; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1952; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1953; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1954; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1955; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1956; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1957; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1958; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1959; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1960; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1961; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1962; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1963; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1964; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1965; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1966; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1967; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1968; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1969; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1970; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1971; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1972; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1973; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1974; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1975; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1976; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1977; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1978; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1979; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1980; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1981; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1982; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1983; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1984; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1985; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1986; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1987; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1988; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1989; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1990; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1991; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1992; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1993; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1994; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1995; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1996; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1997; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1998; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_1999; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2000; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2001; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2002; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2003; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2004; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2005; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2006; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2007; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2008; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2009; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2010; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2011; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2012; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2013; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2014; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2015; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2016; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2017; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2018; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2019; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2020; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2021; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2022; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2023; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2024; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2025; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2026; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2027; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2028; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2029; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2030; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2031; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2032; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2033; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2034; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2035; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2036; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2037; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2038; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2039; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2040; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2041; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2042; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2043; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2044; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2045; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2046; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2047; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2048; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2049; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2050; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2051; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2052; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2053; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2054; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2055; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2056; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2057; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2058; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2059; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2060; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2061; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2062; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2063; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2064; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2065; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2066; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2067; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2068; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2069; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2070; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2071; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2072; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2073; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2074; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2075; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2076; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2077; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2078; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2079; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2080; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2081; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2082; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2083; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2084; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2085; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2086; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2087; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2088; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2089; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2090; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2091; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2092; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2093; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2094; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2095; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2096; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2097; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2098; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2099; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2100; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2101; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2102; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2103; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2104; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2105; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2106; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2107; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2108; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2109; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2110; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2111; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2112; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2113; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2114; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2115; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2116; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2117; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2118; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2119; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2120; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2121; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2122; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2123; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2124; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2125; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2126; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2127; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2128; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2129; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2130; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2131; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2132; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2133; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2134; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2135; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2136; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2137; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2138; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2139; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2140; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2141; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2142; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2143; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2144; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2145; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2146; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2147; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2148; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2149; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2150; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2151; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2152; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2153; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2154; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2155; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2156; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2157; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2158; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2159; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2160; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2161; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2162; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2163; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2164; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2165; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2166; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2167; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2168; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2169; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2170; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2171; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2172; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2173; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2174; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2175; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2176; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2177; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2178; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2179; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2180; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2181; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2182; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2183; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2184; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2185; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2186; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2187; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2188; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2189; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2190; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2191; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2192; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2193; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2194; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2195; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2196; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2197; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2198; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2199; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2200; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2201; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2202; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2203; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2204; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2205; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2206; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2207; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2208; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2209; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2210; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2211; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2212; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2213; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2214; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2215; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2216; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2217; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2218; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2219; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2220; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2221; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2222; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2223; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2224; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2225; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2226; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2227; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2228; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2229; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2230; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2231; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2232; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2233; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2234; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2235; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2236; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2237; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2238; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2239; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2240; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2241; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2242; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2243; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2244; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2245; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2246; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2247; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2248; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2249; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2250; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2251; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2252; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2253; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2254; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2255; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2256; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2257; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2258; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2259; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2260; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2261; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2262; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2263; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2264; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2265; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2266; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2267; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2268; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2269; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2270; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2271; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2272; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2273; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2274; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2275; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2276; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2277; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2278; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2279; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2280; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2281; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2282; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2283; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2284; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2285; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2286; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2287; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2288; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2289; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2290; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2291; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2292; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2293; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2294; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2295; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2296; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2297; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2298; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2299; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2300; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2301; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2302; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2303; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2304; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2305; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2306; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2307; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2308; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2309; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2310; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2311; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2312; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2313; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2314; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2315; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2316; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2317; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2318; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2319; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2320; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2321; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2322; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2323; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2324; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2325; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2326; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2327; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2328; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2329; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2330; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2331; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2332; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2333; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2334; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2335; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2336; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2337; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2338; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2339; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2340; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2341; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2342; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2343; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2344; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2345; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2346; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2347; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2348; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2349; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2350; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2351; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2352; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2353; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2354; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2355; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2356; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2357; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2358; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2359; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2360; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2361; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2362; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2363; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2364; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2365; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2366; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2367; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2368; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2369; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2370; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2371; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2372; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2373; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2374; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2375; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2376; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2377; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2378; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2379; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2380; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2381; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2382; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2383; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2384; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2385; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2386; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2387; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2388; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2389; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2390; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2391; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2392; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2393; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2394; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2395; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2396; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2397; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2398; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2399; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2400; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2401; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2402; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2403; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2404; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2405; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2406; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2407; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2408; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2409; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2410; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2411; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2412; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2413; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2414; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2415; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2416; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2417; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2418; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2419; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2420; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2421; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2422; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2423; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2424; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2425; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2426; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2427; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2428; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2429; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2430; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2431; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2432; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2433; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2434; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2435; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2436; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2437; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2438; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2439; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2440; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2441; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2442; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2443; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2444; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2445; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2446; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2447; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2448; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2449; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2450; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2451; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2452; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2453; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2454; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2455; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2456; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2457; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2458; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2459; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2460; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2461; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2462; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2463; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2464; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2465; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2466; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2467; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2468; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2469; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2470; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2471; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2472; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2473; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2474; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2475; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2476; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2477; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2478; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2479; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2480; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2481; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2482; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2483; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2484; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2485; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2486; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2487; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2488; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2489; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2490; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2491; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2492; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2493; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2494; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2495; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2496; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2497; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2498; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2499; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2500; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2501; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2502; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2503; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2504; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2505; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2506; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2507; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2508; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2509; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2510; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2511; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2512; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2513; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2514; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2515; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2516; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2517; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2518; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2519; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2520; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2521; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2522; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2523; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2524; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2525; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2526; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2527; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2528; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2529; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2530; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2531; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2532; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2533; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2534; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2535; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2536; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2537; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2538; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2539; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2540; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2541; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2542; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2543; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2544; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2545; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2546; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2547; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2548; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2549; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2550; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2551; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2552; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2553; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2554; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2555; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2556; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2557; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2558; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2559; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2560; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2561; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2562; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2563; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2564; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2565; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2566; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2567; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2568; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2569; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2570; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2571; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2572; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2573; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2574; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2575; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2576; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2577; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2578; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2579; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2580; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2581; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2582; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2583; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2584; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2585; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2586; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2587; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2588; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2589; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2590; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2591; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2592; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2593; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2594; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2595; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2596; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2597; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2598; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2599; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2600; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2601; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2602; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2603; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2604; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2605; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2606; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2607; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2608; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2609; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2610; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2611; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2612; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2613; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2614; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2615; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2616; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2617; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2618; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2619; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2620; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2621; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2622; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2623; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2624; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2625; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2626; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2627; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2628; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2629; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2630; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2631; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2632; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2633; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2634; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2635; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2636; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2637; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2638; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2639; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2640; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2641; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2642; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2643; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2644; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2645; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2646; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2647; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2648; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2649; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2650; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2651; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2652; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2653; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2654; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2655; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2656; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2657; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2658; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2659; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2660; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2661; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2662; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2663; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2664; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2665; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2666; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2667; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2668; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2669; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2670; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2671; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2672; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2673; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2674; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2675; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2676; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2677; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2678; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2679; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2680; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2681; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2682; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2683; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2684; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2685; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2686; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2687; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2688; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2689; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2690; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2691; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2692; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2693; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2694; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2695; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2696; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2697; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2698; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2699; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2700; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2701; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2702; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2703; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2704; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2705; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2706; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2707; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2708; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2709; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2710; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2711; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2712; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2713; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2714; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2715; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2716; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2717; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2718; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2719; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2720; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2721; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2722; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2723; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2724; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2725; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2726; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2727; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2728; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2729; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2730; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2731; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2732; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2733; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2734; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2735; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2736; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2737; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2738; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2739; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2740; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2741; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2742; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2743; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2744; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2745; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2746; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2747; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2748; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2749; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2750; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2751; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2752; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2753; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2754; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2755; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2756; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2757; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2758; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2759; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2760; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2761; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2762; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2763; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2764; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2765; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2766; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2767; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2768; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2769; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2770; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2771; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2772; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2773; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2774; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2775; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2776; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2777; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2778; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2779; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2780; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2781; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2782; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2783; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2784; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2785; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2786; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2787; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2788; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2789; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2790; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2791; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2792; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2793; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2794; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2795; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2796; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2797; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2798; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2799; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2800; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2801; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2802; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2803; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2804; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2805; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2806; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2807; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2808; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2809; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2810; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2811; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2812; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2813; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2814; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2815; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2816; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2817; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2818; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2819; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2820; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2821; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2822; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2823; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2824; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2825; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2826; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2827; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2828; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2829; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2830; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2831; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2832; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2833; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2834; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2835; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2836; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2837; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2838; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2839; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2840; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2841; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2842; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2843; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2844; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2845; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2846; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2847; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2848; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2849; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2850; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2851; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2852; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2853; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2854; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2855; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2856; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2857; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2858; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2859; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2860; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2861; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2862; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2863; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2864; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2865; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2866; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2867; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2868; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2869; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2870; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2871; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2872; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2873; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2874; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2875; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2876; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2877; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2878; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2879; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2880; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2881; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2882; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2883; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2884; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2885; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2886; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2887; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2888; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2889; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2890; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2891; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2892; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2893; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2894; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2895; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2896; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2897; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2898; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2899; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2900; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2901; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2902; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2903; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2904; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2905; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2906; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2907; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2908; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2909; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2910; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2911; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2912; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2913; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2914; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2915; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2916; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2917; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2918; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2919; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2920; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2921; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2922; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2923; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2924; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2925; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2926; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2927; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2928; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2929; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2930; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2931; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2932; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2933; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2934; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2935; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2936; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2937; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2938; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2939; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2940; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2941; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2942; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2943; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2944; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2945; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2946; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2947; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2948; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2949; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2950; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2951; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2952; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2953; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2954; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2955; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2956; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2957; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2958; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2959; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2960; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2961; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2962; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2963; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2964; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2965; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2966; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2967; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2968; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2969; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2970; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2971; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2972; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2973; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2974; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2975; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2976; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2977; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2978; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2979; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2980; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2981; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2982; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2983; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2984; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2985; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2986; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2987; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2988; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2989; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2990; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2991; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2992; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2993; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2994; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2995; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2996; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2997; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2998; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_2999; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3000; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3001; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3002; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3003; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3004; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3005; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3006; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3007; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3008; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3009; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3010; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3011; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3012; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3013; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3014; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3015; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3016; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3017; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3018; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3019; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3020; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3021; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3022; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3023; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3024; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3025; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3026; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3027; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3028; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3029; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3030; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3031; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3032; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3033; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3034; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3035; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3036; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3037; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3038; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3039; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3040; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3041; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3042; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3043; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3044; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3045; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3046; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3047; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3048; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3049; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3050; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3051; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3052; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3053; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3054; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3055; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3056; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3057; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3058; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3059; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3060; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3061; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3062; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3063; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3064; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3065; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3066; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3067; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3068; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3069; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3070; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3071; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3072; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3073; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3074; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3075; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3076; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3077; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3078; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3079; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3080; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3081; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3082; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3083; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3084; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3085; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3086; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3087; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3088; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3089; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3090; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3091; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3092; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3093; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3094; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3095; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3096; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3097; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3098; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3099; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3100; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3101; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3102; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3103; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3104; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3105; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3106; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3107; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3108; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3109; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3110; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3111; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3112; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3113; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3114; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3115; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3116; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3117; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3118; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3119; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3120; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3121; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3122; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3123; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3124; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3125; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3126; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3127; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3128; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3129; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3130; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3131; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3132; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3133; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3134; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3135; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3136; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3137; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3138; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3139; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3140; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3141; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3142; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3143; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3144; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3145; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3146; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3147; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3148; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3149; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3150; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3151; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3152; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3153; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3154; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3155; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3156; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3157; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3158; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3159; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3160; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3161; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3162; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3163; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3164; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3165; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3166; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3167; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3168; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3169; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3170; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3171; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3172; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3173; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3174; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3175; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3176; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3177; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3178; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3179; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3180; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3181; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3182; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3183; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3184; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3185; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3186; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3187; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3188; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3189; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3190; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3191; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3192; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3193; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3194; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3195; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3196; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3197; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3198; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3199; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3200; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3201; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3202; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3203; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3204; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3205; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3206; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3207; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3208; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3209; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3210; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3211; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3212; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3213; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3214; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3215; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3216; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3217; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3218; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3219; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3220; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3221; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3222; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3223; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3224; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3225; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3226; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3227; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3228; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3229; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3230; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3231; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3232; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3233; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3234; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3235; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3236; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3237; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3238; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3239; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3240; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3241; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3242; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3243; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3244; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3245; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3246; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3247; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3248; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3249; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3250; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3251; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3252; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3253; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3254; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3255; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3256; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3257; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3258; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3259; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3260; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3261; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3262; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3263; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3264; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3265; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3266; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3267; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3268; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3269; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3270; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3271; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3272; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3273; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3274; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3275; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3276; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3277; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3278; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3279; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3280; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3281; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3282; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3283; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3284; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3285; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3286; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3287; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3288; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3289; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3290; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3291; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3292; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3293; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3294; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3295; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3296; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3297; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3298; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3299; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3300; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3301; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3302; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3303; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3304; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3305; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3306; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3307; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3308; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3309; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3310; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3311; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3312; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3313; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3314; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3315; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3316; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3317; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3318; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3319; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3320; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3321; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3322; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3323; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3324; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3325; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3326; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3327; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3328; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3329; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3330; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3331; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3332; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3333; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3334; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3335; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3336; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3337; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3338; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3339; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3340; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3341; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3342; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3343; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3344; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3345; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3346; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3347; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3348; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3349; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3350; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3351; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3352; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3353; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3354; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3355; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3356; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3357; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3358; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3359; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3360; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3361; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3362; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3363; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3364; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3365; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3366; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3367; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3368; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3369; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3370; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3371; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3372; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3373; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3374; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3375; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3376; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3377; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3378; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3379; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3380; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3381; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3382; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3383; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3384; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3385; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3386; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3387; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3388; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3389; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3390; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3391; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3392; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3393; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3394; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3395; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3396; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3397; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3398; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3399; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3400; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3401; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3402; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3403; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3404; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3405; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3406; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3407; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3408; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3409; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3410; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3411; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3412; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3413; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3414; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3415; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3416; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3417; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3418; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3419; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3420; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3421; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3422; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3423; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3424; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3425; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3426; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3427; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3428; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3429; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3430; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3431; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3432; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3433; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3434; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3435; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3436; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3437; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3438; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3439; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3440; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3441; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3442; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3443; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3444; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3445; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3446; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3447; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3448; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3449; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3450; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3451; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3452; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3453; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3454; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3455; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3456; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3457; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3458; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3459; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3460; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3461; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3462; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3463; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3464; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3465; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3466; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3467; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3468; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3469; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3470; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3471; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3472; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3473; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3474; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3475; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3476; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3477; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3478; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3479; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3480; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3481; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3482; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3483; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3484; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3485; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3486; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3487; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3488; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3489; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3490; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3491; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3492; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3493; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3494; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3495; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3496; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3497; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3498; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3499; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3500; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3501; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3502; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3503; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3504; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3505; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3506; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3507; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3508; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3509; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3510; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3511; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3512; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3513; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3514; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3515; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3516; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3517; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3518; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3519; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3520; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3521; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3522; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3523; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3524; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3525; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3526; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3527; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3528; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3529; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3530; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3531; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3532; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3533; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3534; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3535; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3536; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3537; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3538; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3539; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3540; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3541; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3542; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3543; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3544; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3545; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3546; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3547; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3548; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3549; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3550; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3551; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3552; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3553; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3554; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3555; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3556; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3557; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3558; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3559; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3560; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3561; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3562; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3563; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3564; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3565; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3566; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3567; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3568; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3569; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3570; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3571; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3572; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3573; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3574; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3575; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3576; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3577; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3578; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3579; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3580; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3581; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3582; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3583; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3584; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3585; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3586; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3587; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3588; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3589; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3590; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3591; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3592; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3593; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3594; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3595; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3596; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3597; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3598; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3599; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3600; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3601; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3602; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3603; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3604; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3605; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3606; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3607; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3608; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3609; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3610; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3611; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3612; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3613; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3614; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3615; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3616; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3617; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3618; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3619; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3620; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3621; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3622; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3623; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3624; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3625; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3626; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3627; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3628; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3629; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3630; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3631; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3632; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3633; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3634; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3635; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3636; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3637; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3638; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3639; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3640; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3641; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3642; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3643; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3644; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3645; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3646; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3647; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3648; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3649; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3650; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3651; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3652; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3653; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3654; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3655; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3656; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3657; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3658; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3659; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3660; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3661; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3662; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3663; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3664; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3665; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3666; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3667; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3668; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3669; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3670; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3671; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3672; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3673; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3674; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3675; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3676; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3677; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3678; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3679; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3680; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3681; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3682; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3683; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3684; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3685; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3686; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3687; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3688; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3689; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3690; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3691; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3692; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3693; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3694; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3695; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3696; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3697; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3698; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3699; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3700; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3701; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3702; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3703; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3704; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3705; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3706; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3707; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3708; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3709; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3710; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3711; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3712; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3713; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3714; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3715; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3716; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3717; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3718; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3719; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3720; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3721; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3722; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3723; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3724; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3725; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3726; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3727; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3728; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3729; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3730; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3731; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3732; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3733; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3734; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3735; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3736; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3737; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3738; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3739; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3740; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3741; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3742; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3743; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3744; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3745; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3746; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3747; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3748; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3749; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3750; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3751; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3752; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3753; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3754; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3755; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3756; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3757; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3758; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3759; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3760; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3761; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3762; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3763; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3764; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3765; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3766; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3767; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3768; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3769; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3770; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3771; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3772; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3773; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3774; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3775; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3776; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3777; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3778; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3779; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3780; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3781; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3782; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3783; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3784; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3785; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3786; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3787; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3788; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3789; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3790; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3791; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3792; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3793; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3794; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3795; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3796; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3797; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3798; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3799; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3800; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3801; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3802; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3803; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3804; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3805; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3806; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3807; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3808; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3809; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3810; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3811; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3812; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3813; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3814; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3815; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3816; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3817; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3818; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3819; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3820; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3821; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3822; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3823; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3824; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3825; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3826; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3827; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3828; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3829; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3830; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3831; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3832; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3833; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3834; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3835; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3836; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3837; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3838; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3839; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3840; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3841; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3842; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3843; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3844; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3845; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3846; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3847; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3848; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3849; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3850; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3851; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3852; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3853; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3854; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3855; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3856; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3857; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3858; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3859; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3860; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3861; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3862; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3863; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3864; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3865; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3866; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3867; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3868; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3869; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3870; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3871; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3872; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3873; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3874; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3875; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3876; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3877; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3878; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3879; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3880; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3881; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3882; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3883; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3884; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3885; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3886; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3887; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3888; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3889; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3890; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3891; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3892; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3893; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3894; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3895; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3896; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3897; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3898; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3899; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3900; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3901; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3902; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3903; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3904; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3905; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3906; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3907; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3908; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3909; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3910; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3911; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3912; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3913; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3914; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3915; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3916; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3917; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3918; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3919; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3920; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3921; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3922; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3923; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3924; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3925; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3926; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3927; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3928; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3929; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3930; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3931; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3932; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3933; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3934; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3935; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3936; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3937; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3938; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3939; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3940; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3941; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3942; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3943; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3944; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3945; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3946; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3947; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3948; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3949; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3950; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3951; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3952; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3953; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3954; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3955; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3956; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3957; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3958; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3959; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3960; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3961; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3962; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3963; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3964; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3965; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3966; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3967; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3968; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3969; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3970; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3971; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3972; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3973; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3974; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3975; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3976; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3977; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3978; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3979; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3980; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3981; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3982; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3983; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3984; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3985; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3986; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3987; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3988; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3989; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3990; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3991; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3992; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3993; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3994; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3995; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3996; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3997; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3998; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_3999; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4000; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4001; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4002; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4003; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4004; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4005; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4006; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4007; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4008; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4009; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4010; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4011; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4012; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4013; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4014; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4015; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4016; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4017; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4018; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4019; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4020; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4021; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4022; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4023; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4024; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4025; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4026; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4027; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4028; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4029; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4030; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4031; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4032; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4033; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4034; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4035; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4036; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4037; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4038; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4039; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4040; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4041; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4042; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4043; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4044; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4045; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4046; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4047; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4048; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4049; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4050; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4051; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4052; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4053; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4054; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4055; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4056; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4057; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4058; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4059; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4060; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4061; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4062; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4063; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4064; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4065; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4066; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4067; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4068; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4069; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4070; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4071; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4072; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4073; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4074; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4075; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4076; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4077; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4078; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4079; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4080; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4081; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4082; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4083; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4084; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4085; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4086; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4087; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4088; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4089; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4090; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4091; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4092; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4093; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4094; // @[CSR.scala 31:26]
  reg [31:0] reg_csr_4095; // @[CSR.scala 31:26]
  wire  _csr_addr_T = io_in_id_io_csr_cmd == 3'h4; // @[CSR.scala 40:18]
  wire [31:0] csr_addr = _csr_addr_T ? 32'h342 : io_in_id_io_csr_addr_default; // @[Mux.scala 98:16]
  wire  _csr_wdata_T = io_in_id_io_csr_cmd == 3'h1; // @[CSR.scala 44:18]
  wire  _csr_wdata_T_1 = io_in_id_io_csr_cmd == 3'h2; // @[CSR.scala 45:18]
  wire [31:0] _GEN_1 = 12'h1 == csr_addr[11:0] ? reg_csr_1 : reg_csr_0; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2 = 12'h2 == csr_addr[11:0] ? reg_csr_2 : _GEN_1; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3 = 12'h3 == csr_addr[11:0] ? reg_csr_3 : _GEN_2; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4 = 12'h4 == csr_addr[11:0] ? reg_csr_4 : _GEN_3; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_5 = 12'h5 == csr_addr[11:0] ? reg_csr_5 : _GEN_4; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_6 = 12'h6 == csr_addr[11:0] ? reg_csr_6 : _GEN_5; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_7 = 12'h7 == csr_addr[11:0] ? reg_csr_7 : _GEN_6; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_8 = 12'h8 == csr_addr[11:0] ? reg_csr_8 : _GEN_7; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_9 = 12'h9 == csr_addr[11:0] ? reg_csr_9 : _GEN_8; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_10 = 12'ha == csr_addr[11:0] ? reg_csr_10 : _GEN_9; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_11 = 12'hb == csr_addr[11:0] ? reg_csr_11 : _GEN_10; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_12 = 12'hc == csr_addr[11:0] ? reg_csr_12 : _GEN_11; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_13 = 12'hd == csr_addr[11:0] ? reg_csr_13 : _GEN_12; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_14 = 12'he == csr_addr[11:0] ? reg_csr_14 : _GEN_13; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_15 = 12'hf == csr_addr[11:0] ? reg_csr_15 : _GEN_14; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_16 = 12'h10 == csr_addr[11:0] ? reg_csr_16 : _GEN_15; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_17 = 12'h11 == csr_addr[11:0] ? reg_csr_17 : _GEN_16; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_18 = 12'h12 == csr_addr[11:0] ? reg_csr_18 : _GEN_17; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_19 = 12'h13 == csr_addr[11:0] ? reg_csr_19 : _GEN_18; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_20 = 12'h14 == csr_addr[11:0] ? reg_csr_20 : _GEN_19; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_21 = 12'h15 == csr_addr[11:0] ? reg_csr_21 : _GEN_20; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_22 = 12'h16 == csr_addr[11:0] ? reg_csr_22 : _GEN_21; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_23 = 12'h17 == csr_addr[11:0] ? reg_csr_23 : _GEN_22; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_24 = 12'h18 == csr_addr[11:0] ? reg_csr_24 : _GEN_23; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_25 = 12'h19 == csr_addr[11:0] ? reg_csr_25 : _GEN_24; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_26 = 12'h1a == csr_addr[11:0] ? reg_csr_26 : _GEN_25; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_27 = 12'h1b == csr_addr[11:0] ? reg_csr_27 : _GEN_26; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_28 = 12'h1c == csr_addr[11:0] ? reg_csr_28 : _GEN_27; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_29 = 12'h1d == csr_addr[11:0] ? reg_csr_29 : _GEN_28; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_30 = 12'h1e == csr_addr[11:0] ? reg_csr_30 : _GEN_29; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_31 = 12'h1f == csr_addr[11:0] ? reg_csr_31 : _GEN_30; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_32 = 12'h20 == csr_addr[11:0] ? reg_csr_32 : _GEN_31; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_33 = 12'h21 == csr_addr[11:0] ? reg_csr_33 : _GEN_32; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_34 = 12'h22 == csr_addr[11:0] ? reg_csr_34 : _GEN_33; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_35 = 12'h23 == csr_addr[11:0] ? reg_csr_35 : _GEN_34; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_36 = 12'h24 == csr_addr[11:0] ? reg_csr_36 : _GEN_35; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_37 = 12'h25 == csr_addr[11:0] ? reg_csr_37 : _GEN_36; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_38 = 12'h26 == csr_addr[11:0] ? reg_csr_38 : _GEN_37; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_39 = 12'h27 == csr_addr[11:0] ? reg_csr_39 : _GEN_38; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_40 = 12'h28 == csr_addr[11:0] ? reg_csr_40 : _GEN_39; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_41 = 12'h29 == csr_addr[11:0] ? reg_csr_41 : _GEN_40; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_42 = 12'h2a == csr_addr[11:0] ? reg_csr_42 : _GEN_41; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_43 = 12'h2b == csr_addr[11:0] ? reg_csr_43 : _GEN_42; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_44 = 12'h2c == csr_addr[11:0] ? reg_csr_44 : _GEN_43; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_45 = 12'h2d == csr_addr[11:0] ? reg_csr_45 : _GEN_44; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_46 = 12'h2e == csr_addr[11:0] ? reg_csr_46 : _GEN_45; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_47 = 12'h2f == csr_addr[11:0] ? reg_csr_47 : _GEN_46; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_48 = 12'h30 == csr_addr[11:0] ? reg_csr_48 : _GEN_47; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_49 = 12'h31 == csr_addr[11:0] ? reg_csr_49 : _GEN_48; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_50 = 12'h32 == csr_addr[11:0] ? reg_csr_50 : _GEN_49; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_51 = 12'h33 == csr_addr[11:0] ? reg_csr_51 : _GEN_50; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_52 = 12'h34 == csr_addr[11:0] ? reg_csr_52 : _GEN_51; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_53 = 12'h35 == csr_addr[11:0] ? reg_csr_53 : _GEN_52; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_54 = 12'h36 == csr_addr[11:0] ? reg_csr_54 : _GEN_53; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_55 = 12'h37 == csr_addr[11:0] ? reg_csr_55 : _GEN_54; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_56 = 12'h38 == csr_addr[11:0] ? reg_csr_56 : _GEN_55; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_57 = 12'h39 == csr_addr[11:0] ? reg_csr_57 : _GEN_56; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_58 = 12'h3a == csr_addr[11:0] ? reg_csr_58 : _GEN_57; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_59 = 12'h3b == csr_addr[11:0] ? reg_csr_59 : _GEN_58; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_60 = 12'h3c == csr_addr[11:0] ? reg_csr_60 : _GEN_59; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_61 = 12'h3d == csr_addr[11:0] ? reg_csr_61 : _GEN_60; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_62 = 12'h3e == csr_addr[11:0] ? reg_csr_62 : _GEN_61; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_63 = 12'h3f == csr_addr[11:0] ? reg_csr_63 : _GEN_62; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_64 = 12'h40 == csr_addr[11:0] ? reg_csr_64 : _GEN_63; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_65 = 12'h41 == csr_addr[11:0] ? reg_csr_65 : _GEN_64; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_66 = 12'h42 == csr_addr[11:0] ? reg_csr_66 : _GEN_65; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_67 = 12'h43 == csr_addr[11:0] ? reg_csr_67 : _GEN_66; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_68 = 12'h44 == csr_addr[11:0] ? reg_csr_68 : _GEN_67; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_69 = 12'h45 == csr_addr[11:0] ? reg_csr_69 : _GEN_68; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_70 = 12'h46 == csr_addr[11:0] ? reg_csr_70 : _GEN_69; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_71 = 12'h47 == csr_addr[11:0] ? reg_csr_71 : _GEN_70; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_72 = 12'h48 == csr_addr[11:0] ? reg_csr_72 : _GEN_71; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_73 = 12'h49 == csr_addr[11:0] ? reg_csr_73 : _GEN_72; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_74 = 12'h4a == csr_addr[11:0] ? reg_csr_74 : _GEN_73; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_75 = 12'h4b == csr_addr[11:0] ? reg_csr_75 : _GEN_74; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_76 = 12'h4c == csr_addr[11:0] ? reg_csr_76 : _GEN_75; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_77 = 12'h4d == csr_addr[11:0] ? reg_csr_77 : _GEN_76; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_78 = 12'h4e == csr_addr[11:0] ? reg_csr_78 : _GEN_77; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_79 = 12'h4f == csr_addr[11:0] ? reg_csr_79 : _GEN_78; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_80 = 12'h50 == csr_addr[11:0] ? reg_csr_80 : _GEN_79; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_81 = 12'h51 == csr_addr[11:0] ? reg_csr_81 : _GEN_80; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_82 = 12'h52 == csr_addr[11:0] ? reg_csr_82 : _GEN_81; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_83 = 12'h53 == csr_addr[11:0] ? reg_csr_83 : _GEN_82; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_84 = 12'h54 == csr_addr[11:0] ? reg_csr_84 : _GEN_83; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_85 = 12'h55 == csr_addr[11:0] ? reg_csr_85 : _GEN_84; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_86 = 12'h56 == csr_addr[11:0] ? reg_csr_86 : _GEN_85; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_87 = 12'h57 == csr_addr[11:0] ? reg_csr_87 : _GEN_86; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_88 = 12'h58 == csr_addr[11:0] ? reg_csr_88 : _GEN_87; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_89 = 12'h59 == csr_addr[11:0] ? reg_csr_89 : _GEN_88; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_90 = 12'h5a == csr_addr[11:0] ? reg_csr_90 : _GEN_89; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_91 = 12'h5b == csr_addr[11:0] ? reg_csr_91 : _GEN_90; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_92 = 12'h5c == csr_addr[11:0] ? reg_csr_92 : _GEN_91; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_93 = 12'h5d == csr_addr[11:0] ? reg_csr_93 : _GEN_92; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_94 = 12'h5e == csr_addr[11:0] ? reg_csr_94 : _GEN_93; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_95 = 12'h5f == csr_addr[11:0] ? reg_csr_95 : _GEN_94; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_96 = 12'h60 == csr_addr[11:0] ? reg_csr_96 : _GEN_95; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_97 = 12'h61 == csr_addr[11:0] ? reg_csr_97 : _GEN_96; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_98 = 12'h62 == csr_addr[11:0] ? reg_csr_98 : _GEN_97; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_99 = 12'h63 == csr_addr[11:0] ? reg_csr_99 : _GEN_98; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_100 = 12'h64 == csr_addr[11:0] ? reg_csr_100 : _GEN_99; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_101 = 12'h65 == csr_addr[11:0] ? reg_csr_101 : _GEN_100; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_102 = 12'h66 == csr_addr[11:0] ? reg_csr_102 : _GEN_101; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_103 = 12'h67 == csr_addr[11:0] ? reg_csr_103 : _GEN_102; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_104 = 12'h68 == csr_addr[11:0] ? reg_csr_104 : _GEN_103; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_105 = 12'h69 == csr_addr[11:0] ? reg_csr_105 : _GEN_104; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_106 = 12'h6a == csr_addr[11:0] ? reg_csr_106 : _GEN_105; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_107 = 12'h6b == csr_addr[11:0] ? reg_csr_107 : _GEN_106; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_108 = 12'h6c == csr_addr[11:0] ? reg_csr_108 : _GEN_107; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_109 = 12'h6d == csr_addr[11:0] ? reg_csr_109 : _GEN_108; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_110 = 12'h6e == csr_addr[11:0] ? reg_csr_110 : _GEN_109; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_111 = 12'h6f == csr_addr[11:0] ? reg_csr_111 : _GEN_110; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_112 = 12'h70 == csr_addr[11:0] ? reg_csr_112 : _GEN_111; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_113 = 12'h71 == csr_addr[11:0] ? reg_csr_113 : _GEN_112; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_114 = 12'h72 == csr_addr[11:0] ? reg_csr_114 : _GEN_113; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_115 = 12'h73 == csr_addr[11:0] ? reg_csr_115 : _GEN_114; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_116 = 12'h74 == csr_addr[11:0] ? reg_csr_116 : _GEN_115; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_117 = 12'h75 == csr_addr[11:0] ? reg_csr_117 : _GEN_116; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_118 = 12'h76 == csr_addr[11:0] ? reg_csr_118 : _GEN_117; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_119 = 12'h77 == csr_addr[11:0] ? reg_csr_119 : _GEN_118; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_120 = 12'h78 == csr_addr[11:0] ? reg_csr_120 : _GEN_119; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_121 = 12'h79 == csr_addr[11:0] ? reg_csr_121 : _GEN_120; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_122 = 12'h7a == csr_addr[11:0] ? reg_csr_122 : _GEN_121; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_123 = 12'h7b == csr_addr[11:0] ? reg_csr_123 : _GEN_122; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_124 = 12'h7c == csr_addr[11:0] ? reg_csr_124 : _GEN_123; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_125 = 12'h7d == csr_addr[11:0] ? reg_csr_125 : _GEN_124; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_126 = 12'h7e == csr_addr[11:0] ? reg_csr_126 : _GEN_125; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_127 = 12'h7f == csr_addr[11:0] ? reg_csr_127 : _GEN_126; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_128 = 12'h80 == csr_addr[11:0] ? reg_csr_128 : _GEN_127; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_129 = 12'h81 == csr_addr[11:0] ? reg_csr_129 : _GEN_128; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_130 = 12'h82 == csr_addr[11:0] ? reg_csr_130 : _GEN_129; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_131 = 12'h83 == csr_addr[11:0] ? reg_csr_131 : _GEN_130; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_132 = 12'h84 == csr_addr[11:0] ? reg_csr_132 : _GEN_131; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_133 = 12'h85 == csr_addr[11:0] ? reg_csr_133 : _GEN_132; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_134 = 12'h86 == csr_addr[11:0] ? reg_csr_134 : _GEN_133; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_135 = 12'h87 == csr_addr[11:0] ? reg_csr_135 : _GEN_134; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_136 = 12'h88 == csr_addr[11:0] ? reg_csr_136 : _GEN_135; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_137 = 12'h89 == csr_addr[11:0] ? reg_csr_137 : _GEN_136; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_138 = 12'h8a == csr_addr[11:0] ? reg_csr_138 : _GEN_137; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_139 = 12'h8b == csr_addr[11:0] ? reg_csr_139 : _GEN_138; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_140 = 12'h8c == csr_addr[11:0] ? reg_csr_140 : _GEN_139; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_141 = 12'h8d == csr_addr[11:0] ? reg_csr_141 : _GEN_140; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_142 = 12'h8e == csr_addr[11:0] ? reg_csr_142 : _GEN_141; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_143 = 12'h8f == csr_addr[11:0] ? reg_csr_143 : _GEN_142; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_144 = 12'h90 == csr_addr[11:0] ? reg_csr_144 : _GEN_143; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_145 = 12'h91 == csr_addr[11:0] ? reg_csr_145 : _GEN_144; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_146 = 12'h92 == csr_addr[11:0] ? reg_csr_146 : _GEN_145; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_147 = 12'h93 == csr_addr[11:0] ? reg_csr_147 : _GEN_146; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_148 = 12'h94 == csr_addr[11:0] ? reg_csr_148 : _GEN_147; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_149 = 12'h95 == csr_addr[11:0] ? reg_csr_149 : _GEN_148; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_150 = 12'h96 == csr_addr[11:0] ? reg_csr_150 : _GEN_149; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_151 = 12'h97 == csr_addr[11:0] ? reg_csr_151 : _GEN_150; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_152 = 12'h98 == csr_addr[11:0] ? reg_csr_152 : _GEN_151; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_153 = 12'h99 == csr_addr[11:0] ? reg_csr_153 : _GEN_152; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_154 = 12'h9a == csr_addr[11:0] ? reg_csr_154 : _GEN_153; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_155 = 12'h9b == csr_addr[11:0] ? reg_csr_155 : _GEN_154; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_156 = 12'h9c == csr_addr[11:0] ? reg_csr_156 : _GEN_155; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_157 = 12'h9d == csr_addr[11:0] ? reg_csr_157 : _GEN_156; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_158 = 12'h9e == csr_addr[11:0] ? reg_csr_158 : _GEN_157; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_159 = 12'h9f == csr_addr[11:0] ? reg_csr_159 : _GEN_158; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_160 = 12'ha0 == csr_addr[11:0] ? reg_csr_160 : _GEN_159; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_161 = 12'ha1 == csr_addr[11:0] ? reg_csr_161 : _GEN_160; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_162 = 12'ha2 == csr_addr[11:0] ? reg_csr_162 : _GEN_161; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_163 = 12'ha3 == csr_addr[11:0] ? reg_csr_163 : _GEN_162; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_164 = 12'ha4 == csr_addr[11:0] ? reg_csr_164 : _GEN_163; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_165 = 12'ha5 == csr_addr[11:0] ? reg_csr_165 : _GEN_164; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_166 = 12'ha6 == csr_addr[11:0] ? reg_csr_166 : _GEN_165; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_167 = 12'ha7 == csr_addr[11:0] ? reg_csr_167 : _GEN_166; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_168 = 12'ha8 == csr_addr[11:0] ? reg_csr_168 : _GEN_167; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_169 = 12'ha9 == csr_addr[11:0] ? reg_csr_169 : _GEN_168; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_170 = 12'haa == csr_addr[11:0] ? reg_csr_170 : _GEN_169; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_171 = 12'hab == csr_addr[11:0] ? reg_csr_171 : _GEN_170; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_172 = 12'hac == csr_addr[11:0] ? reg_csr_172 : _GEN_171; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_173 = 12'had == csr_addr[11:0] ? reg_csr_173 : _GEN_172; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_174 = 12'hae == csr_addr[11:0] ? reg_csr_174 : _GEN_173; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_175 = 12'haf == csr_addr[11:0] ? reg_csr_175 : _GEN_174; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_176 = 12'hb0 == csr_addr[11:0] ? reg_csr_176 : _GEN_175; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_177 = 12'hb1 == csr_addr[11:0] ? reg_csr_177 : _GEN_176; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_178 = 12'hb2 == csr_addr[11:0] ? reg_csr_178 : _GEN_177; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_179 = 12'hb3 == csr_addr[11:0] ? reg_csr_179 : _GEN_178; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_180 = 12'hb4 == csr_addr[11:0] ? reg_csr_180 : _GEN_179; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_181 = 12'hb5 == csr_addr[11:0] ? reg_csr_181 : _GEN_180; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_182 = 12'hb6 == csr_addr[11:0] ? reg_csr_182 : _GEN_181; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_183 = 12'hb7 == csr_addr[11:0] ? reg_csr_183 : _GEN_182; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_184 = 12'hb8 == csr_addr[11:0] ? reg_csr_184 : _GEN_183; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_185 = 12'hb9 == csr_addr[11:0] ? reg_csr_185 : _GEN_184; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_186 = 12'hba == csr_addr[11:0] ? reg_csr_186 : _GEN_185; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_187 = 12'hbb == csr_addr[11:0] ? reg_csr_187 : _GEN_186; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_188 = 12'hbc == csr_addr[11:0] ? reg_csr_188 : _GEN_187; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_189 = 12'hbd == csr_addr[11:0] ? reg_csr_189 : _GEN_188; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_190 = 12'hbe == csr_addr[11:0] ? reg_csr_190 : _GEN_189; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_191 = 12'hbf == csr_addr[11:0] ? reg_csr_191 : _GEN_190; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_192 = 12'hc0 == csr_addr[11:0] ? reg_csr_192 : _GEN_191; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_193 = 12'hc1 == csr_addr[11:0] ? reg_csr_193 : _GEN_192; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_194 = 12'hc2 == csr_addr[11:0] ? reg_csr_194 : _GEN_193; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_195 = 12'hc3 == csr_addr[11:0] ? reg_csr_195 : _GEN_194; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_196 = 12'hc4 == csr_addr[11:0] ? reg_csr_196 : _GEN_195; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_197 = 12'hc5 == csr_addr[11:0] ? reg_csr_197 : _GEN_196; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_198 = 12'hc6 == csr_addr[11:0] ? reg_csr_198 : _GEN_197; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_199 = 12'hc7 == csr_addr[11:0] ? reg_csr_199 : _GEN_198; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_200 = 12'hc8 == csr_addr[11:0] ? reg_csr_200 : _GEN_199; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_201 = 12'hc9 == csr_addr[11:0] ? reg_csr_201 : _GEN_200; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_202 = 12'hca == csr_addr[11:0] ? reg_csr_202 : _GEN_201; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_203 = 12'hcb == csr_addr[11:0] ? reg_csr_203 : _GEN_202; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_204 = 12'hcc == csr_addr[11:0] ? reg_csr_204 : _GEN_203; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_205 = 12'hcd == csr_addr[11:0] ? reg_csr_205 : _GEN_204; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_206 = 12'hce == csr_addr[11:0] ? reg_csr_206 : _GEN_205; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_207 = 12'hcf == csr_addr[11:0] ? reg_csr_207 : _GEN_206; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_208 = 12'hd0 == csr_addr[11:0] ? reg_csr_208 : _GEN_207; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_209 = 12'hd1 == csr_addr[11:0] ? reg_csr_209 : _GEN_208; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_210 = 12'hd2 == csr_addr[11:0] ? reg_csr_210 : _GEN_209; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_211 = 12'hd3 == csr_addr[11:0] ? reg_csr_211 : _GEN_210; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_212 = 12'hd4 == csr_addr[11:0] ? reg_csr_212 : _GEN_211; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_213 = 12'hd5 == csr_addr[11:0] ? reg_csr_213 : _GEN_212; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_214 = 12'hd6 == csr_addr[11:0] ? reg_csr_214 : _GEN_213; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_215 = 12'hd7 == csr_addr[11:0] ? reg_csr_215 : _GEN_214; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_216 = 12'hd8 == csr_addr[11:0] ? reg_csr_216 : _GEN_215; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_217 = 12'hd9 == csr_addr[11:0] ? reg_csr_217 : _GEN_216; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_218 = 12'hda == csr_addr[11:0] ? reg_csr_218 : _GEN_217; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_219 = 12'hdb == csr_addr[11:0] ? reg_csr_219 : _GEN_218; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_220 = 12'hdc == csr_addr[11:0] ? reg_csr_220 : _GEN_219; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_221 = 12'hdd == csr_addr[11:0] ? reg_csr_221 : _GEN_220; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_222 = 12'hde == csr_addr[11:0] ? reg_csr_222 : _GEN_221; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_223 = 12'hdf == csr_addr[11:0] ? reg_csr_223 : _GEN_222; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_224 = 12'he0 == csr_addr[11:0] ? reg_csr_224 : _GEN_223; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_225 = 12'he1 == csr_addr[11:0] ? reg_csr_225 : _GEN_224; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_226 = 12'he2 == csr_addr[11:0] ? reg_csr_226 : _GEN_225; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_227 = 12'he3 == csr_addr[11:0] ? reg_csr_227 : _GEN_226; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_228 = 12'he4 == csr_addr[11:0] ? reg_csr_228 : _GEN_227; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_229 = 12'he5 == csr_addr[11:0] ? reg_csr_229 : _GEN_228; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_230 = 12'he6 == csr_addr[11:0] ? reg_csr_230 : _GEN_229; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_231 = 12'he7 == csr_addr[11:0] ? reg_csr_231 : _GEN_230; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_232 = 12'he8 == csr_addr[11:0] ? reg_csr_232 : _GEN_231; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_233 = 12'he9 == csr_addr[11:0] ? reg_csr_233 : _GEN_232; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_234 = 12'hea == csr_addr[11:0] ? reg_csr_234 : _GEN_233; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_235 = 12'heb == csr_addr[11:0] ? reg_csr_235 : _GEN_234; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_236 = 12'hec == csr_addr[11:0] ? reg_csr_236 : _GEN_235; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_237 = 12'hed == csr_addr[11:0] ? reg_csr_237 : _GEN_236; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_238 = 12'hee == csr_addr[11:0] ? reg_csr_238 : _GEN_237; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_239 = 12'hef == csr_addr[11:0] ? reg_csr_239 : _GEN_238; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_240 = 12'hf0 == csr_addr[11:0] ? reg_csr_240 : _GEN_239; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_241 = 12'hf1 == csr_addr[11:0] ? reg_csr_241 : _GEN_240; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_242 = 12'hf2 == csr_addr[11:0] ? reg_csr_242 : _GEN_241; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_243 = 12'hf3 == csr_addr[11:0] ? reg_csr_243 : _GEN_242; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_244 = 12'hf4 == csr_addr[11:0] ? reg_csr_244 : _GEN_243; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_245 = 12'hf5 == csr_addr[11:0] ? reg_csr_245 : _GEN_244; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_246 = 12'hf6 == csr_addr[11:0] ? reg_csr_246 : _GEN_245; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_247 = 12'hf7 == csr_addr[11:0] ? reg_csr_247 : _GEN_246; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_248 = 12'hf8 == csr_addr[11:0] ? reg_csr_248 : _GEN_247; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_249 = 12'hf9 == csr_addr[11:0] ? reg_csr_249 : _GEN_248; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_250 = 12'hfa == csr_addr[11:0] ? reg_csr_250 : _GEN_249; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_251 = 12'hfb == csr_addr[11:0] ? reg_csr_251 : _GEN_250; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_252 = 12'hfc == csr_addr[11:0] ? reg_csr_252 : _GEN_251; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_253 = 12'hfd == csr_addr[11:0] ? reg_csr_253 : _GEN_252; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_254 = 12'hfe == csr_addr[11:0] ? reg_csr_254 : _GEN_253; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_255 = 12'hff == csr_addr[11:0] ? reg_csr_255 : _GEN_254; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_256 = 12'h100 == csr_addr[11:0] ? reg_csr_256 : _GEN_255; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_257 = 12'h101 == csr_addr[11:0] ? reg_csr_257 : _GEN_256; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_258 = 12'h102 == csr_addr[11:0] ? reg_csr_258 : _GEN_257; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_259 = 12'h103 == csr_addr[11:0] ? reg_csr_259 : _GEN_258; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_260 = 12'h104 == csr_addr[11:0] ? reg_csr_260 : _GEN_259; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_261 = 12'h105 == csr_addr[11:0] ? reg_csr_261 : _GEN_260; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_262 = 12'h106 == csr_addr[11:0] ? reg_csr_262 : _GEN_261; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_263 = 12'h107 == csr_addr[11:0] ? reg_csr_263 : _GEN_262; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_264 = 12'h108 == csr_addr[11:0] ? reg_csr_264 : _GEN_263; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_265 = 12'h109 == csr_addr[11:0] ? reg_csr_265 : _GEN_264; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_266 = 12'h10a == csr_addr[11:0] ? reg_csr_266 : _GEN_265; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_267 = 12'h10b == csr_addr[11:0] ? reg_csr_267 : _GEN_266; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_268 = 12'h10c == csr_addr[11:0] ? reg_csr_268 : _GEN_267; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_269 = 12'h10d == csr_addr[11:0] ? reg_csr_269 : _GEN_268; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_270 = 12'h10e == csr_addr[11:0] ? reg_csr_270 : _GEN_269; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_271 = 12'h10f == csr_addr[11:0] ? reg_csr_271 : _GEN_270; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_272 = 12'h110 == csr_addr[11:0] ? reg_csr_272 : _GEN_271; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_273 = 12'h111 == csr_addr[11:0] ? reg_csr_273 : _GEN_272; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_274 = 12'h112 == csr_addr[11:0] ? reg_csr_274 : _GEN_273; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_275 = 12'h113 == csr_addr[11:0] ? reg_csr_275 : _GEN_274; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_276 = 12'h114 == csr_addr[11:0] ? reg_csr_276 : _GEN_275; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_277 = 12'h115 == csr_addr[11:0] ? reg_csr_277 : _GEN_276; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_278 = 12'h116 == csr_addr[11:0] ? reg_csr_278 : _GEN_277; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_279 = 12'h117 == csr_addr[11:0] ? reg_csr_279 : _GEN_278; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_280 = 12'h118 == csr_addr[11:0] ? reg_csr_280 : _GEN_279; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_281 = 12'h119 == csr_addr[11:0] ? reg_csr_281 : _GEN_280; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_282 = 12'h11a == csr_addr[11:0] ? reg_csr_282 : _GEN_281; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_283 = 12'h11b == csr_addr[11:0] ? reg_csr_283 : _GEN_282; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_284 = 12'h11c == csr_addr[11:0] ? reg_csr_284 : _GEN_283; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_285 = 12'h11d == csr_addr[11:0] ? reg_csr_285 : _GEN_284; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_286 = 12'h11e == csr_addr[11:0] ? reg_csr_286 : _GEN_285; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_287 = 12'h11f == csr_addr[11:0] ? reg_csr_287 : _GEN_286; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_288 = 12'h120 == csr_addr[11:0] ? reg_csr_288 : _GEN_287; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_289 = 12'h121 == csr_addr[11:0] ? reg_csr_289 : _GEN_288; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_290 = 12'h122 == csr_addr[11:0] ? reg_csr_290 : _GEN_289; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_291 = 12'h123 == csr_addr[11:0] ? reg_csr_291 : _GEN_290; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_292 = 12'h124 == csr_addr[11:0] ? reg_csr_292 : _GEN_291; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_293 = 12'h125 == csr_addr[11:0] ? reg_csr_293 : _GEN_292; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_294 = 12'h126 == csr_addr[11:0] ? reg_csr_294 : _GEN_293; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_295 = 12'h127 == csr_addr[11:0] ? reg_csr_295 : _GEN_294; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_296 = 12'h128 == csr_addr[11:0] ? reg_csr_296 : _GEN_295; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_297 = 12'h129 == csr_addr[11:0] ? reg_csr_297 : _GEN_296; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_298 = 12'h12a == csr_addr[11:0] ? reg_csr_298 : _GEN_297; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_299 = 12'h12b == csr_addr[11:0] ? reg_csr_299 : _GEN_298; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_300 = 12'h12c == csr_addr[11:0] ? reg_csr_300 : _GEN_299; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_301 = 12'h12d == csr_addr[11:0] ? reg_csr_301 : _GEN_300; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_302 = 12'h12e == csr_addr[11:0] ? reg_csr_302 : _GEN_301; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_303 = 12'h12f == csr_addr[11:0] ? reg_csr_303 : _GEN_302; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_304 = 12'h130 == csr_addr[11:0] ? reg_csr_304 : _GEN_303; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_305 = 12'h131 == csr_addr[11:0] ? reg_csr_305 : _GEN_304; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_306 = 12'h132 == csr_addr[11:0] ? reg_csr_306 : _GEN_305; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_307 = 12'h133 == csr_addr[11:0] ? reg_csr_307 : _GEN_306; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_308 = 12'h134 == csr_addr[11:0] ? reg_csr_308 : _GEN_307; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_309 = 12'h135 == csr_addr[11:0] ? reg_csr_309 : _GEN_308; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_310 = 12'h136 == csr_addr[11:0] ? reg_csr_310 : _GEN_309; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_311 = 12'h137 == csr_addr[11:0] ? reg_csr_311 : _GEN_310; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_312 = 12'h138 == csr_addr[11:0] ? reg_csr_312 : _GEN_311; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_313 = 12'h139 == csr_addr[11:0] ? reg_csr_313 : _GEN_312; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_314 = 12'h13a == csr_addr[11:0] ? reg_csr_314 : _GEN_313; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_315 = 12'h13b == csr_addr[11:0] ? reg_csr_315 : _GEN_314; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_316 = 12'h13c == csr_addr[11:0] ? reg_csr_316 : _GEN_315; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_317 = 12'h13d == csr_addr[11:0] ? reg_csr_317 : _GEN_316; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_318 = 12'h13e == csr_addr[11:0] ? reg_csr_318 : _GEN_317; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_319 = 12'h13f == csr_addr[11:0] ? reg_csr_319 : _GEN_318; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_320 = 12'h140 == csr_addr[11:0] ? reg_csr_320 : _GEN_319; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_321 = 12'h141 == csr_addr[11:0] ? reg_csr_321 : _GEN_320; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_322 = 12'h142 == csr_addr[11:0] ? reg_csr_322 : _GEN_321; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_323 = 12'h143 == csr_addr[11:0] ? reg_csr_323 : _GEN_322; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_324 = 12'h144 == csr_addr[11:0] ? reg_csr_324 : _GEN_323; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_325 = 12'h145 == csr_addr[11:0] ? reg_csr_325 : _GEN_324; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_326 = 12'h146 == csr_addr[11:0] ? reg_csr_326 : _GEN_325; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_327 = 12'h147 == csr_addr[11:0] ? reg_csr_327 : _GEN_326; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_328 = 12'h148 == csr_addr[11:0] ? reg_csr_328 : _GEN_327; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_329 = 12'h149 == csr_addr[11:0] ? reg_csr_329 : _GEN_328; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_330 = 12'h14a == csr_addr[11:0] ? reg_csr_330 : _GEN_329; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_331 = 12'h14b == csr_addr[11:0] ? reg_csr_331 : _GEN_330; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_332 = 12'h14c == csr_addr[11:0] ? reg_csr_332 : _GEN_331; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_333 = 12'h14d == csr_addr[11:0] ? reg_csr_333 : _GEN_332; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_334 = 12'h14e == csr_addr[11:0] ? reg_csr_334 : _GEN_333; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_335 = 12'h14f == csr_addr[11:0] ? reg_csr_335 : _GEN_334; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_336 = 12'h150 == csr_addr[11:0] ? reg_csr_336 : _GEN_335; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_337 = 12'h151 == csr_addr[11:0] ? reg_csr_337 : _GEN_336; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_338 = 12'h152 == csr_addr[11:0] ? reg_csr_338 : _GEN_337; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_339 = 12'h153 == csr_addr[11:0] ? reg_csr_339 : _GEN_338; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_340 = 12'h154 == csr_addr[11:0] ? reg_csr_340 : _GEN_339; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_341 = 12'h155 == csr_addr[11:0] ? reg_csr_341 : _GEN_340; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_342 = 12'h156 == csr_addr[11:0] ? reg_csr_342 : _GEN_341; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_343 = 12'h157 == csr_addr[11:0] ? reg_csr_343 : _GEN_342; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_344 = 12'h158 == csr_addr[11:0] ? reg_csr_344 : _GEN_343; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_345 = 12'h159 == csr_addr[11:0] ? reg_csr_345 : _GEN_344; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_346 = 12'h15a == csr_addr[11:0] ? reg_csr_346 : _GEN_345; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_347 = 12'h15b == csr_addr[11:0] ? reg_csr_347 : _GEN_346; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_348 = 12'h15c == csr_addr[11:0] ? reg_csr_348 : _GEN_347; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_349 = 12'h15d == csr_addr[11:0] ? reg_csr_349 : _GEN_348; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_350 = 12'h15e == csr_addr[11:0] ? reg_csr_350 : _GEN_349; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_351 = 12'h15f == csr_addr[11:0] ? reg_csr_351 : _GEN_350; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_352 = 12'h160 == csr_addr[11:0] ? reg_csr_352 : _GEN_351; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_353 = 12'h161 == csr_addr[11:0] ? reg_csr_353 : _GEN_352; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_354 = 12'h162 == csr_addr[11:0] ? reg_csr_354 : _GEN_353; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_355 = 12'h163 == csr_addr[11:0] ? reg_csr_355 : _GEN_354; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_356 = 12'h164 == csr_addr[11:0] ? reg_csr_356 : _GEN_355; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_357 = 12'h165 == csr_addr[11:0] ? reg_csr_357 : _GEN_356; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_358 = 12'h166 == csr_addr[11:0] ? reg_csr_358 : _GEN_357; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_359 = 12'h167 == csr_addr[11:0] ? reg_csr_359 : _GEN_358; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_360 = 12'h168 == csr_addr[11:0] ? reg_csr_360 : _GEN_359; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_361 = 12'h169 == csr_addr[11:0] ? reg_csr_361 : _GEN_360; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_362 = 12'h16a == csr_addr[11:0] ? reg_csr_362 : _GEN_361; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_363 = 12'h16b == csr_addr[11:0] ? reg_csr_363 : _GEN_362; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_364 = 12'h16c == csr_addr[11:0] ? reg_csr_364 : _GEN_363; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_365 = 12'h16d == csr_addr[11:0] ? reg_csr_365 : _GEN_364; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_366 = 12'h16e == csr_addr[11:0] ? reg_csr_366 : _GEN_365; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_367 = 12'h16f == csr_addr[11:0] ? reg_csr_367 : _GEN_366; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_368 = 12'h170 == csr_addr[11:0] ? reg_csr_368 : _GEN_367; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_369 = 12'h171 == csr_addr[11:0] ? reg_csr_369 : _GEN_368; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_370 = 12'h172 == csr_addr[11:0] ? reg_csr_370 : _GEN_369; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_371 = 12'h173 == csr_addr[11:0] ? reg_csr_371 : _GEN_370; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_372 = 12'h174 == csr_addr[11:0] ? reg_csr_372 : _GEN_371; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_373 = 12'h175 == csr_addr[11:0] ? reg_csr_373 : _GEN_372; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_374 = 12'h176 == csr_addr[11:0] ? reg_csr_374 : _GEN_373; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_375 = 12'h177 == csr_addr[11:0] ? reg_csr_375 : _GEN_374; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_376 = 12'h178 == csr_addr[11:0] ? reg_csr_376 : _GEN_375; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_377 = 12'h179 == csr_addr[11:0] ? reg_csr_377 : _GEN_376; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_378 = 12'h17a == csr_addr[11:0] ? reg_csr_378 : _GEN_377; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_379 = 12'h17b == csr_addr[11:0] ? reg_csr_379 : _GEN_378; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_380 = 12'h17c == csr_addr[11:0] ? reg_csr_380 : _GEN_379; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_381 = 12'h17d == csr_addr[11:0] ? reg_csr_381 : _GEN_380; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_382 = 12'h17e == csr_addr[11:0] ? reg_csr_382 : _GEN_381; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_383 = 12'h17f == csr_addr[11:0] ? reg_csr_383 : _GEN_382; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_384 = 12'h180 == csr_addr[11:0] ? reg_csr_384 : _GEN_383; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_385 = 12'h181 == csr_addr[11:0] ? reg_csr_385 : _GEN_384; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_386 = 12'h182 == csr_addr[11:0] ? reg_csr_386 : _GEN_385; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_387 = 12'h183 == csr_addr[11:0] ? reg_csr_387 : _GEN_386; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_388 = 12'h184 == csr_addr[11:0] ? reg_csr_388 : _GEN_387; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_389 = 12'h185 == csr_addr[11:0] ? reg_csr_389 : _GEN_388; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_390 = 12'h186 == csr_addr[11:0] ? reg_csr_390 : _GEN_389; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_391 = 12'h187 == csr_addr[11:0] ? reg_csr_391 : _GEN_390; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_392 = 12'h188 == csr_addr[11:0] ? reg_csr_392 : _GEN_391; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_393 = 12'h189 == csr_addr[11:0] ? reg_csr_393 : _GEN_392; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_394 = 12'h18a == csr_addr[11:0] ? reg_csr_394 : _GEN_393; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_395 = 12'h18b == csr_addr[11:0] ? reg_csr_395 : _GEN_394; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_396 = 12'h18c == csr_addr[11:0] ? reg_csr_396 : _GEN_395; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_397 = 12'h18d == csr_addr[11:0] ? reg_csr_397 : _GEN_396; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_398 = 12'h18e == csr_addr[11:0] ? reg_csr_398 : _GEN_397; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_399 = 12'h18f == csr_addr[11:0] ? reg_csr_399 : _GEN_398; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_400 = 12'h190 == csr_addr[11:0] ? reg_csr_400 : _GEN_399; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_401 = 12'h191 == csr_addr[11:0] ? reg_csr_401 : _GEN_400; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_402 = 12'h192 == csr_addr[11:0] ? reg_csr_402 : _GEN_401; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_403 = 12'h193 == csr_addr[11:0] ? reg_csr_403 : _GEN_402; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_404 = 12'h194 == csr_addr[11:0] ? reg_csr_404 : _GEN_403; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_405 = 12'h195 == csr_addr[11:0] ? reg_csr_405 : _GEN_404; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_406 = 12'h196 == csr_addr[11:0] ? reg_csr_406 : _GEN_405; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_407 = 12'h197 == csr_addr[11:0] ? reg_csr_407 : _GEN_406; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_408 = 12'h198 == csr_addr[11:0] ? reg_csr_408 : _GEN_407; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_409 = 12'h199 == csr_addr[11:0] ? reg_csr_409 : _GEN_408; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_410 = 12'h19a == csr_addr[11:0] ? reg_csr_410 : _GEN_409; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_411 = 12'h19b == csr_addr[11:0] ? reg_csr_411 : _GEN_410; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_412 = 12'h19c == csr_addr[11:0] ? reg_csr_412 : _GEN_411; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_413 = 12'h19d == csr_addr[11:0] ? reg_csr_413 : _GEN_412; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_414 = 12'h19e == csr_addr[11:0] ? reg_csr_414 : _GEN_413; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_415 = 12'h19f == csr_addr[11:0] ? reg_csr_415 : _GEN_414; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_416 = 12'h1a0 == csr_addr[11:0] ? reg_csr_416 : _GEN_415; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_417 = 12'h1a1 == csr_addr[11:0] ? reg_csr_417 : _GEN_416; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_418 = 12'h1a2 == csr_addr[11:0] ? reg_csr_418 : _GEN_417; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_419 = 12'h1a3 == csr_addr[11:0] ? reg_csr_419 : _GEN_418; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_420 = 12'h1a4 == csr_addr[11:0] ? reg_csr_420 : _GEN_419; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_421 = 12'h1a5 == csr_addr[11:0] ? reg_csr_421 : _GEN_420; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_422 = 12'h1a6 == csr_addr[11:0] ? reg_csr_422 : _GEN_421; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_423 = 12'h1a7 == csr_addr[11:0] ? reg_csr_423 : _GEN_422; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_424 = 12'h1a8 == csr_addr[11:0] ? reg_csr_424 : _GEN_423; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_425 = 12'h1a9 == csr_addr[11:0] ? reg_csr_425 : _GEN_424; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_426 = 12'h1aa == csr_addr[11:0] ? reg_csr_426 : _GEN_425; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_427 = 12'h1ab == csr_addr[11:0] ? reg_csr_427 : _GEN_426; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_428 = 12'h1ac == csr_addr[11:0] ? reg_csr_428 : _GEN_427; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_429 = 12'h1ad == csr_addr[11:0] ? reg_csr_429 : _GEN_428; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_430 = 12'h1ae == csr_addr[11:0] ? reg_csr_430 : _GEN_429; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_431 = 12'h1af == csr_addr[11:0] ? reg_csr_431 : _GEN_430; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_432 = 12'h1b0 == csr_addr[11:0] ? reg_csr_432 : _GEN_431; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_433 = 12'h1b1 == csr_addr[11:0] ? reg_csr_433 : _GEN_432; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_434 = 12'h1b2 == csr_addr[11:0] ? reg_csr_434 : _GEN_433; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_435 = 12'h1b3 == csr_addr[11:0] ? reg_csr_435 : _GEN_434; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_436 = 12'h1b4 == csr_addr[11:0] ? reg_csr_436 : _GEN_435; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_437 = 12'h1b5 == csr_addr[11:0] ? reg_csr_437 : _GEN_436; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_438 = 12'h1b6 == csr_addr[11:0] ? reg_csr_438 : _GEN_437; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_439 = 12'h1b7 == csr_addr[11:0] ? reg_csr_439 : _GEN_438; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_440 = 12'h1b8 == csr_addr[11:0] ? reg_csr_440 : _GEN_439; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_441 = 12'h1b9 == csr_addr[11:0] ? reg_csr_441 : _GEN_440; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_442 = 12'h1ba == csr_addr[11:0] ? reg_csr_442 : _GEN_441; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_443 = 12'h1bb == csr_addr[11:0] ? reg_csr_443 : _GEN_442; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_444 = 12'h1bc == csr_addr[11:0] ? reg_csr_444 : _GEN_443; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_445 = 12'h1bd == csr_addr[11:0] ? reg_csr_445 : _GEN_444; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_446 = 12'h1be == csr_addr[11:0] ? reg_csr_446 : _GEN_445; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_447 = 12'h1bf == csr_addr[11:0] ? reg_csr_447 : _GEN_446; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_448 = 12'h1c0 == csr_addr[11:0] ? reg_csr_448 : _GEN_447; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_449 = 12'h1c1 == csr_addr[11:0] ? reg_csr_449 : _GEN_448; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_450 = 12'h1c2 == csr_addr[11:0] ? reg_csr_450 : _GEN_449; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_451 = 12'h1c3 == csr_addr[11:0] ? reg_csr_451 : _GEN_450; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_452 = 12'h1c4 == csr_addr[11:0] ? reg_csr_452 : _GEN_451; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_453 = 12'h1c5 == csr_addr[11:0] ? reg_csr_453 : _GEN_452; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_454 = 12'h1c6 == csr_addr[11:0] ? reg_csr_454 : _GEN_453; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_455 = 12'h1c7 == csr_addr[11:0] ? reg_csr_455 : _GEN_454; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_456 = 12'h1c8 == csr_addr[11:0] ? reg_csr_456 : _GEN_455; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_457 = 12'h1c9 == csr_addr[11:0] ? reg_csr_457 : _GEN_456; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_458 = 12'h1ca == csr_addr[11:0] ? reg_csr_458 : _GEN_457; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_459 = 12'h1cb == csr_addr[11:0] ? reg_csr_459 : _GEN_458; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_460 = 12'h1cc == csr_addr[11:0] ? reg_csr_460 : _GEN_459; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_461 = 12'h1cd == csr_addr[11:0] ? reg_csr_461 : _GEN_460; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_462 = 12'h1ce == csr_addr[11:0] ? reg_csr_462 : _GEN_461; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_463 = 12'h1cf == csr_addr[11:0] ? reg_csr_463 : _GEN_462; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_464 = 12'h1d0 == csr_addr[11:0] ? reg_csr_464 : _GEN_463; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_465 = 12'h1d1 == csr_addr[11:0] ? reg_csr_465 : _GEN_464; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_466 = 12'h1d2 == csr_addr[11:0] ? reg_csr_466 : _GEN_465; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_467 = 12'h1d3 == csr_addr[11:0] ? reg_csr_467 : _GEN_466; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_468 = 12'h1d4 == csr_addr[11:0] ? reg_csr_468 : _GEN_467; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_469 = 12'h1d5 == csr_addr[11:0] ? reg_csr_469 : _GEN_468; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_470 = 12'h1d6 == csr_addr[11:0] ? reg_csr_470 : _GEN_469; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_471 = 12'h1d7 == csr_addr[11:0] ? reg_csr_471 : _GEN_470; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_472 = 12'h1d8 == csr_addr[11:0] ? reg_csr_472 : _GEN_471; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_473 = 12'h1d9 == csr_addr[11:0] ? reg_csr_473 : _GEN_472; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_474 = 12'h1da == csr_addr[11:0] ? reg_csr_474 : _GEN_473; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_475 = 12'h1db == csr_addr[11:0] ? reg_csr_475 : _GEN_474; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_476 = 12'h1dc == csr_addr[11:0] ? reg_csr_476 : _GEN_475; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_477 = 12'h1dd == csr_addr[11:0] ? reg_csr_477 : _GEN_476; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_478 = 12'h1de == csr_addr[11:0] ? reg_csr_478 : _GEN_477; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_479 = 12'h1df == csr_addr[11:0] ? reg_csr_479 : _GEN_478; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_480 = 12'h1e0 == csr_addr[11:0] ? reg_csr_480 : _GEN_479; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_481 = 12'h1e1 == csr_addr[11:0] ? reg_csr_481 : _GEN_480; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_482 = 12'h1e2 == csr_addr[11:0] ? reg_csr_482 : _GEN_481; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_483 = 12'h1e3 == csr_addr[11:0] ? reg_csr_483 : _GEN_482; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_484 = 12'h1e4 == csr_addr[11:0] ? reg_csr_484 : _GEN_483; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_485 = 12'h1e5 == csr_addr[11:0] ? reg_csr_485 : _GEN_484; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_486 = 12'h1e6 == csr_addr[11:0] ? reg_csr_486 : _GEN_485; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_487 = 12'h1e7 == csr_addr[11:0] ? reg_csr_487 : _GEN_486; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_488 = 12'h1e8 == csr_addr[11:0] ? reg_csr_488 : _GEN_487; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_489 = 12'h1e9 == csr_addr[11:0] ? reg_csr_489 : _GEN_488; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_490 = 12'h1ea == csr_addr[11:0] ? reg_csr_490 : _GEN_489; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_491 = 12'h1eb == csr_addr[11:0] ? reg_csr_491 : _GEN_490; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_492 = 12'h1ec == csr_addr[11:0] ? reg_csr_492 : _GEN_491; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_493 = 12'h1ed == csr_addr[11:0] ? reg_csr_493 : _GEN_492; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_494 = 12'h1ee == csr_addr[11:0] ? reg_csr_494 : _GEN_493; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_495 = 12'h1ef == csr_addr[11:0] ? reg_csr_495 : _GEN_494; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_496 = 12'h1f0 == csr_addr[11:0] ? reg_csr_496 : _GEN_495; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_497 = 12'h1f1 == csr_addr[11:0] ? reg_csr_497 : _GEN_496; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_498 = 12'h1f2 == csr_addr[11:0] ? reg_csr_498 : _GEN_497; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_499 = 12'h1f3 == csr_addr[11:0] ? reg_csr_499 : _GEN_498; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_500 = 12'h1f4 == csr_addr[11:0] ? reg_csr_500 : _GEN_499; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_501 = 12'h1f5 == csr_addr[11:0] ? reg_csr_501 : _GEN_500; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_502 = 12'h1f6 == csr_addr[11:0] ? reg_csr_502 : _GEN_501; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_503 = 12'h1f7 == csr_addr[11:0] ? reg_csr_503 : _GEN_502; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_504 = 12'h1f8 == csr_addr[11:0] ? reg_csr_504 : _GEN_503; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_505 = 12'h1f9 == csr_addr[11:0] ? reg_csr_505 : _GEN_504; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_506 = 12'h1fa == csr_addr[11:0] ? reg_csr_506 : _GEN_505; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_507 = 12'h1fb == csr_addr[11:0] ? reg_csr_507 : _GEN_506; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_508 = 12'h1fc == csr_addr[11:0] ? reg_csr_508 : _GEN_507; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_509 = 12'h1fd == csr_addr[11:0] ? reg_csr_509 : _GEN_508; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_510 = 12'h1fe == csr_addr[11:0] ? reg_csr_510 : _GEN_509; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_511 = 12'h1ff == csr_addr[11:0] ? reg_csr_511 : _GEN_510; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_512 = 12'h200 == csr_addr[11:0] ? reg_csr_512 : _GEN_511; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_513 = 12'h201 == csr_addr[11:0] ? reg_csr_513 : _GEN_512; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_514 = 12'h202 == csr_addr[11:0] ? reg_csr_514 : _GEN_513; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_515 = 12'h203 == csr_addr[11:0] ? reg_csr_515 : _GEN_514; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_516 = 12'h204 == csr_addr[11:0] ? reg_csr_516 : _GEN_515; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_517 = 12'h205 == csr_addr[11:0] ? reg_csr_517 : _GEN_516; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_518 = 12'h206 == csr_addr[11:0] ? reg_csr_518 : _GEN_517; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_519 = 12'h207 == csr_addr[11:0] ? reg_csr_519 : _GEN_518; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_520 = 12'h208 == csr_addr[11:0] ? reg_csr_520 : _GEN_519; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_521 = 12'h209 == csr_addr[11:0] ? reg_csr_521 : _GEN_520; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_522 = 12'h20a == csr_addr[11:0] ? reg_csr_522 : _GEN_521; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_523 = 12'h20b == csr_addr[11:0] ? reg_csr_523 : _GEN_522; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_524 = 12'h20c == csr_addr[11:0] ? reg_csr_524 : _GEN_523; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_525 = 12'h20d == csr_addr[11:0] ? reg_csr_525 : _GEN_524; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_526 = 12'h20e == csr_addr[11:0] ? reg_csr_526 : _GEN_525; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_527 = 12'h20f == csr_addr[11:0] ? reg_csr_527 : _GEN_526; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_528 = 12'h210 == csr_addr[11:0] ? reg_csr_528 : _GEN_527; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_529 = 12'h211 == csr_addr[11:0] ? reg_csr_529 : _GEN_528; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_530 = 12'h212 == csr_addr[11:0] ? reg_csr_530 : _GEN_529; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_531 = 12'h213 == csr_addr[11:0] ? reg_csr_531 : _GEN_530; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_532 = 12'h214 == csr_addr[11:0] ? reg_csr_532 : _GEN_531; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_533 = 12'h215 == csr_addr[11:0] ? reg_csr_533 : _GEN_532; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_534 = 12'h216 == csr_addr[11:0] ? reg_csr_534 : _GEN_533; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_535 = 12'h217 == csr_addr[11:0] ? reg_csr_535 : _GEN_534; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_536 = 12'h218 == csr_addr[11:0] ? reg_csr_536 : _GEN_535; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_537 = 12'h219 == csr_addr[11:0] ? reg_csr_537 : _GEN_536; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_538 = 12'h21a == csr_addr[11:0] ? reg_csr_538 : _GEN_537; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_539 = 12'h21b == csr_addr[11:0] ? reg_csr_539 : _GEN_538; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_540 = 12'h21c == csr_addr[11:0] ? reg_csr_540 : _GEN_539; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_541 = 12'h21d == csr_addr[11:0] ? reg_csr_541 : _GEN_540; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_542 = 12'h21e == csr_addr[11:0] ? reg_csr_542 : _GEN_541; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_543 = 12'h21f == csr_addr[11:0] ? reg_csr_543 : _GEN_542; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_544 = 12'h220 == csr_addr[11:0] ? reg_csr_544 : _GEN_543; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_545 = 12'h221 == csr_addr[11:0] ? reg_csr_545 : _GEN_544; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_546 = 12'h222 == csr_addr[11:0] ? reg_csr_546 : _GEN_545; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_547 = 12'h223 == csr_addr[11:0] ? reg_csr_547 : _GEN_546; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_548 = 12'h224 == csr_addr[11:0] ? reg_csr_548 : _GEN_547; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_549 = 12'h225 == csr_addr[11:0] ? reg_csr_549 : _GEN_548; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_550 = 12'h226 == csr_addr[11:0] ? reg_csr_550 : _GEN_549; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_551 = 12'h227 == csr_addr[11:0] ? reg_csr_551 : _GEN_550; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_552 = 12'h228 == csr_addr[11:0] ? reg_csr_552 : _GEN_551; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_553 = 12'h229 == csr_addr[11:0] ? reg_csr_553 : _GEN_552; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_554 = 12'h22a == csr_addr[11:0] ? reg_csr_554 : _GEN_553; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_555 = 12'h22b == csr_addr[11:0] ? reg_csr_555 : _GEN_554; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_556 = 12'h22c == csr_addr[11:0] ? reg_csr_556 : _GEN_555; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_557 = 12'h22d == csr_addr[11:0] ? reg_csr_557 : _GEN_556; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_558 = 12'h22e == csr_addr[11:0] ? reg_csr_558 : _GEN_557; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_559 = 12'h22f == csr_addr[11:0] ? reg_csr_559 : _GEN_558; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_560 = 12'h230 == csr_addr[11:0] ? reg_csr_560 : _GEN_559; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_561 = 12'h231 == csr_addr[11:0] ? reg_csr_561 : _GEN_560; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_562 = 12'h232 == csr_addr[11:0] ? reg_csr_562 : _GEN_561; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_563 = 12'h233 == csr_addr[11:0] ? reg_csr_563 : _GEN_562; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_564 = 12'h234 == csr_addr[11:0] ? reg_csr_564 : _GEN_563; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_565 = 12'h235 == csr_addr[11:0] ? reg_csr_565 : _GEN_564; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_566 = 12'h236 == csr_addr[11:0] ? reg_csr_566 : _GEN_565; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_567 = 12'h237 == csr_addr[11:0] ? reg_csr_567 : _GEN_566; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_568 = 12'h238 == csr_addr[11:0] ? reg_csr_568 : _GEN_567; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_569 = 12'h239 == csr_addr[11:0] ? reg_csr_569 : _GEN_568; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_570 = 12'h23a == csr_addr[11:0] ? reg_csr_570 : _GEN_569; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_571 = 12'h23b == csr_addr[11:0] ? reg_csr_571 : _GEN_570; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_572 = 12'h23c == csr_addr[11:0] ? reg_csr_572 : _GEN_571; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_573 = 12'h23d == csr_addr[11:0] ? reg_csr_573 : _GEN_572; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_574 = 12'h23e == csr_addr[11:0] ? reg_csr_574 : _GEN_573; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_575 = 12'h23f == csr_addr[11:0] ? reg_csr_575 : _GEN_574; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_576 = 12'h240 == csr_addr[11:0] ? reg_csr_576 : _GEN_575; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_577 = 12'h241 == csr_addr[11:0] ? reg_csr_577 : _GEN_576; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_578 = 12'h242 == csr_addr[11:0] ? reg_csr_578 : _GEN_577; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_579 = 12'h243 == csr_addr[11:0] ? reg_csr_579 : _GEN_578; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_580 = 12'h244 == csr_addr[11:0] ? reg_csr_580 : _GEN_579; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_581 = 12'h245 == csr_addr[11:0] ? reg_csr_581 : _GEN_580; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_582 = 12'h246 == csr_addr[11:0] ? reg_csr_582 : _GEN_581; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_583 = 12'h247 == csr_addr[11:0] ? reg_csr_583 : _GEN_582; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_584 = 12'h248 == csr_addr[11:0] ? reg_csr_584 : _GEN_583; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_585 = 12'h249 == csr_addr[11:0] ? reg_csr_585 : _GEN_584; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_586 = 12'h24a == csr_addr[11:0] ? reg_csr_586 : _GEN_585; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_587 = 12'h24b == csr_addr[11:0] ? reg_csr_587 : _GEN_586; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_588 = 12'h24c == csr_addr[11:0] ? reg_csr_588 : _GEN_587; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_589 = 12'h24d == csr_addr[11:0] ? reg_csr_589 : _GEN_588; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_590 = 12'h24e == csr_addr[11:0] ? reg_csr_590 : _GEN_589; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_591 = 12'h24f == csr_addr[11:0] ? reg_csr_591 : _GEN_590; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_592 = 12'h250 == csr_addr[11:0] ? reg_csr_592 : _GEN_591; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_593 = 12'h251 == csr_addr[11:0] ? reg_csr_593 : _GEN_592; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_594 = 12'h252 == csr_addr[11:0] ? reg_csr_594 : _GEN_593; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_595 = 12'h253 == csr_addr[11:0] ? reg_csr_595 : _GEN_594; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_596 = 12'h254 == csr_addr[11:0] ? reg_csr_596 : _GEN_595; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_597 = 12'h255 == csr_addr[11:0] ? reg_csr_597 : _GEN_596; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_598 = 12'h256 == csr_addr[11:0] ? reg_csr_598 : _GEN_597; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_599 = 12'h257 == csr_addr[11:0] ? reg_csr_599 : _GEN_598; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_600 = 12'h258 == csr_addr[11:0] ? reg_csr_600 : _GEN_599; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_601 = 12'h259 == csr_addr[11:0] ? reg_csr_601 : _GEN_600; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_602 = 12'h25a == csr_addr[11:0] ? reg_csr_602 : _GEN_601; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_603 = 12'h25b == csr_addr[11:0] ? reg_csr_603 : _GEN_602; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_604 = 12'h25c == csr_addr[11:0] ? reg_csr_604 : _GEN_603; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_605 = 12'h25d == csr_addr[11:0] ? reg_csr_605 : _GEN_604; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_606 = 12'h25e == csr_addr[11:0] ? reg_csr_606 : _GEN_605; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_607 = 12'h25f == csr_addr[11:0] ? reg_csr_607 : _GEN_606; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_608 = 12'h260 == csr_addr[11:0] ? reg_csr_608 : _GEN_607; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_609 = 12'h261 == csr_addr[11:0] ? reg_csr_609 : _GEN_608; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_610 = 12'h262 == csr_addr[11:0] ? reg_csr_610 : _GEN_609; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_611 = 12'h263 == csr_addr[11:0] ? reg_csr_611 : _GEN_610; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_612 = 12'h264 == csr_addr[11:0] ? reg_csr_612 : _GEN_611; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_613 = 12'h265 == csr_addr[11:0] ? reg_csr_613 : _GEN_612; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_614 = 12'h266 == csr_addr[11:0] ? reg_csr_614 : _GEN_613; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_615 = 12'h267 == csr_addr[11:0] ? reg_csr_615 : _GEN_614; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_616 = 12'h268 == csr_addr[11:0] ? reg_csr_616 : _GEN_615; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_617 = 12'h269 == csr_addr[11:0] ? reg_csr_617 : _GEN_616; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_618 = 12'h26a == csr_addr[11:0] ? reg_csr_618 : _GEN_617; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_619 = 12'h26b == csr_addr[11:0] ? reg_csr_619 : _GEN_618; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_620 = 12'h26c == csr_addr[11:0] ? reg_csr_620 : _GEN_619; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_621 = 12'h26d == csr_addr[11:0] ? reg_csr_621 : _GEN_620; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_622 = 12'h26e == csr_addr[11:0] ? reg_csr_622 : _GEN_621; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_623 = 12'h26f == csr_addr[11:0] ? reg_csr_623 : _GEN_622; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_624 = 12'h270 == csr_addr[11:0] ? reg_csr_624 : _GEN_623; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_625 = 12'h271 == csr_addr[11:0] ? reg_csr_625 : _GEN_624; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_626 = 12'h272 == csr_addr[11:0] ? reg_csr_626 : _GEN_625; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_627 = 12'h273 == csr_addr[11:0] ? reg_csr_627 : _GEN_626; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_628 = 12'h274 == csr_addr[11:0] ? reg_csr_628 : _GEN_627; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_629 = 12'h275 == csr_addr[11:0] ? reg_csr_629 : _GEN_628; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_630 = 12'h276 == csr_addr[11:0] ? reg_csr_630 : _GEN_629; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_631 = 12'h277 == csr_addr[11:0] ? reg_csr_631 : _GEN_630; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_632 = 12'h278 == csr_addr[11:0] ? reg_csr_632 : _GEN_631; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_633 = 12'h279 == csr_addr[11:0] ? reg_csr_633 : _GEN_632; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_634 = 12'h27a == csr_addr[11:0] ? reg_csr_634 : _GEN_633; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_635 = 12'h27b == csr_addr[11:0] ? reg_csr_635 : _GEN_634; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_636 = 12'h27c == csr_addr[11:0] ? reg_csr_636 : _GEN_635; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_637 = 12'h27d == csr_addr[11:0] ? reg_csr_637 : _GEN_636; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_638 = 12'h27e == csr_addr[11:0] ? reg_csr_638 : _GEN_637; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_639 = 12'h27f == csr_addr[11:0] ? reg_csr_639 : _GEN_638; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_640 = 12'h280 == csr_addr[11:0] ? reg_csr_640 : _GEN_639; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_641 = 12'h281 == csr_addr[11:0] ? reg_csr_641 : _GEN_640; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_642 = 12'h282 == csr_addr[11:0] ? reg_csr_642 : _GEN_641; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_643 = 12'h283 == csr_addr[11:0] ? reg_csr_643 : _GEN_642; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_644 = 12'h284 == csr_addr[11:0] ? reg_csr_644 : _GEN_643; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_645 = 12'h285 == csr_addr[11:0] ? reg_csr_645 : _GEN_644; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_646 = 12'h286 == csr_addr[11:0] ? reg_csr_646 : _GEN_645; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_647 = 12'h287 == csr_addr[11:0] ? reg_csr_647 : _GEN_646; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_648 = 12'h288 == csr_addr[11:0] ? reg_csr_648 : _GEN_647; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_649 = 12'h289 == csr_addr[11:0] ? reg_csr_649 : _GEN_648; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_650 = 12'h28a == csr_addr[11:0] ? reg_csr_650 : _GEN_649; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_651 = 12'h28b == csr_addr[11:0] ? reg_csr_651 : _GEN_650; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_652 = 12'h28c == csr_addr[11:0] ? reg_csr_652 : _GEN_651; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_653 = 12'h28d == csr_addr[11:0] ? reg_csr_653 : _GEN_652; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_654 = 12'h28e == csr_addr[11:0] ? reg_csr_654 : _GEN_653; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_655 = 12'h28f == csr_addr[11:0] ? reg_csr_655 : _GEN_654; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_656 = 12'h290 == csr_addr[11:0] ? reg_csr_656 : _GEN_655; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_657 = 12'h291 == csr_addr[11:0] ? reg_csr_657 : _GEN_656; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_658 = 12'h292 == csr_addr[11:0] ? reg_csr_658 : _GEN_657; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_659 = 12'h293 == csr_addr[11:0] ? reg_csr_659 : _GEN_658; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_660 = 12'h294 == csr_addr[11:0] ? reg_csr_660 : _GEN_659; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_661 = 12'h295 == csr_addr[11:0] ? reg_csr_661 : _GEN_660; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_662 = 12'h296 == csr_addr[11:0] ? reg_csr_662 : _GEN_661; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_663 = 12'h297 == csr_addr[11:0] ? reg_csr_663 : _GEN_662; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_664 = 12'h298 == csr_addr[11:0] ? reg_csr_664 : _GEN_663; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_665 = 12'h299 == csr_addr[11:0] ? reg_csr_665 : _GEN_664; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_666 = 12'h29a == csr_addr[11:0] ? reg_csr_666 : _GEN_665; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_667 = 12'h29b == csr_addr[11:0] ? reg_csr_667 : _GEN_666; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_668 = 12'h29c == csr_addr[11:0] ? reg_csr_668 : _GEN_667; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_669 = 12'h29d == csr_addr[11:0] ? reg_csr_669 : _GEN_668; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_670 = 12'h29e == csr_addr[11:0] ? reg_csr_670 : _GEN_669; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_671 = 12'h29f == csr_addr[11:0] ? reg_csr_671 : _GEN_670; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_672 = 12'h2a0 == csr_addr[11:0] ? reg_csr_672 : _GEN_671; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_673 = 12'h2a1 == csr_addr[11:0] ? reg_csr_673 : _GEN_672; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_674 = 12'h2a2 == csr_addr[11:0] ? reg_csr_674 : _GEN_673; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_675 = 12'h2a3 == csr_addr[11:0] ? reg_csr_675 : _GEN_674; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_676 = 12'h2a4 == csr_addr[11:0] ? reg_csr_676 : _GEN_675; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_677 = 12'h2a5 == csr_addr[11:0] ? reg_csr_677 : _GEN_676; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_678 = 12'h2a6 == csr_addr[11:0] ? reg_csr_678 : _GEN_677; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_679 = 12'h2a7 == csr_addr[11:0] ? reg_csr_679 : _GEN_678; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_680 = 12'h2a8 == csr_addr[11:0] ? reg_csr_680 : _GEN_679; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_681 = 12'h2a9 == csr_addr[11:0] ? reg_csr_681 : _GEN_680; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_682 = 12'h2aa == csr_addr[11:0] ? reg_csr_682 : _GEN_681; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_683 = 12'h2ab == csr_addr[11:0] ? reg_csr_683 : _GEN_682; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_684 = 12'h2ac == csr_addr[11:0] ? reg_csr_684 : _GEN_683; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_685 = 12'h2ad == csr_addr[11:0] ? reg_csr_685 : _GEN_684; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_686 = 12'h2ae == csr_addr[11:0] ? reg_csr_686 : _GEN_685; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_687 = 12'h2af == csr_addr[11:0] ? reg_csr_687 : _GEN_686; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_688 = 12'h2b0 == csr_addr[11:0] ? reg_csr_688 : _GEN_687; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_689 = 12'h2b1 == csr_addr[11:0] ? reg_csr_689 : _GEN_688; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_690 = 12'h2b2 == csr_addr[11:0] ? reg_csr_690 : _GEN_689; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_691 = 12'h2b3 == csr_addr[11:0] ? reg_csr_691 : _GEN_690; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_692 = 12'h2b4 == csr_addr[11:0] ? reg_csr_692 : _GEN_691; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_693 = 12'h2b5 == csr_addr[11:0] ? reg_csr_693 : _GEN_692; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_694 = 12'h2b6 == csr_addr[11:0] ? reg_csr_694 : _GEN_693; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_695 = 12'h2b7 == csr_addr[11:0] ? reg_csr_695 : _GEN_694; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_696 = 12'h2b8 == csr_addr[11:0] ? reg_csr_696 : _GEN_695; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_697 = 12'h2b9 == csr_addr[11:0] ? reg_csr_697 : _GEN_696; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_698 = 12'h2ba == csr_addr[11:0] ? reg_csr_698 : _GEN_697; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_699 = 12'h2bb == csr_addr[11:0] ? reg_csr_699 : _GEN_698; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_700 = 12'h2bc == csr_addr[11:0] ? reg_csr_700 : _GEN_699; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_701 = 12'h2bd == csr_addr[11:0] ? reg_csr_701 : _GEN_700; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_702 = 12'h2be == csr_addr[11:0] ? reg_csr_702 : _GEN_701; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_703 = 12'h2bf == csr_addr[11:0] ? reg_csr_703 : _GEN_702; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_704 = 12'h2c0 == csr_addr[11:0] ? reg_csr_704 : _GEN_703; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_705 = 12'h2c1 == csr_addr[11:0] ? reg_csr_705 : _GEN_704; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_706 = 12'h2c2 == csr_addr[11:0] ? reg_csr_706 : _GEN_705; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_707 = 12'h2c3 == csr_addr[11:0] ? reg_csr_707 : _GEN_706; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_708 = 12'h2c4 == csr_addr[11:0] ? reg_csr_708 : _GEN_707; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_709 = 12'h2c5 == csr_addr[11:0] ? reg_csr_709 : _GEN_708; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_710 = 12'h2c6 == csr_addr[11:0] ? reg_csr_710 : _GEN_709; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_711 = 12'h2c7 == csr_addr[11:0] ? reg_csr_711 : _GEN_710; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_712 = 12'h2c8 == csr_addr[11:0] ? reg_csr_712 : _GEN_711; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_713 = 12'h2c9 == csr_addr[11:0] ? reg_csr_713 : _GEN_712; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_714 = 12'h2ca == csr_addr[11:0] ? reg_csr_714 : _GEN_713; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_715 = 12'h2cb == csr_addr[11:0] ? reg_csr_715 : _GEN_714; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_716 = 12'h2cc == csr_addr[11:0] ? reg_csr_716 : _GEN_715; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_717 = 12'h2cd == csr_addr[11:0] ? reg_csr_717 : _GEN_716; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_718 = 12'h2ce == csr_addr[11:0] ? reg_csr_718 : _GEN_717; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_719 = 12'h2cf == csr_addr[11:0] ? reg_csr_719 : _GEN_718; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_720 = 12'h2d0 == csr_addr[11:0] ? reg_csr_720 : _GEN_719; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_721 = 12'h2d1 == csr_addr[11:0] ? reg_csr_721 : _GEN_720; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_722 = 12'h2d2 == csr_addr[11:0] ? reg_csr_722 : _GEN_721; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_723 = 12'h2d3 == csr_addr[11:0] ? reg_csr_723 : _GEN_722; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_724 = 12'h2d4 == csr_addr[11:0] ? reg_csr_724 : _GEN_723; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_725 = 12'h2d5 == csr_addr[11:0] ? reg_csr_725 : _GEN_724; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_726 = 12'h2d6 == csr_addr[11:0] ? reg_csr_726 : _GEN_725; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_727 = 12'h2d7 == csr_addr[11:0] ? reg_csr_727 : _GEN_726; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_728 = 12'h2d8 == csr_addr[11:0] ? reg_csr_728 : _GEN_727; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_729 = 12'h2d9 == csr_addr[11:0] ? reg_csr_729 : _GEN_728; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_730 = 12'h2da == csr_addr[11:0] ? reg_csr_730 : _GEN_729; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_731 = 12'h2db == csr_addr[11:0] ? reg_csr_731 : _GEN_730; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_732 = 12'h2dc == csr_addr[11:0] ? reg_csr_732 : _GEN_731; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_733 = 12'h2dd == csr_addr[11:0] ? reg_csr_733 : _GEN_732; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_734 = 12'h2de == csr_addr[11:0] ? reg_csr_734 : _GEN_733; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_735 = 12'h2df == csr_addr[11:0] ? reg_csr_735 : _GEN_734; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_736 = 12'h2e0 == csr_addr[11:0] ? reg_csr_736 : _GEN_735; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_737 = 12'h2e1 == csr_addr[11:0] ? reg_csr_737 : _GEN_736; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_738 = 12'h2e2 == csr_addr[11:0] ? reg_csr_738 : _GEN_737; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_739 = 12'h2e3 == csr_addr[11:0] ? reg_csr_739 : _GEN_738; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_740 = 12'h2e4 == csr_addr[11:0] ? reg_csr_740 : _GEN_739; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_741 = 12'h2e5 == csr_addr[11:0] ? reg_csr_741 : _GEN_740; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_742 = 12'h2e6 == csr_addr[11:0] ? reg_csr_742 : _GEN_741; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_743 = 12'h2e7 == csr_addr[11:0] ? reg_csr_743 : _GEN_742; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_744 = 12'h2e8 == csr_addr[11:0] ? reg_csr_744 : _GEN_743; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_745 = 12'h2e9 == csr_addr[11:0] ? reg_csr_745 : _GEN_744; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_746 = 12'h2ea == csr_addr[11:0] ? reg_csr_746 : _GEN_745; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_747 = 12'h2eb == csr_addr[11:0] ? reg_csr_747 : _GEN_746; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_748 = 12'h2ec == csr_addr[11:0] ? reg_csr_748 : _GEN_747; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_749 = 12'h2ed == csr_addr[11:0] ? reg_csr_749 : _GEN_748; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_750 = 12'h2ee == csr_addr[11:0] ? reg_csr_750 : _GEN_749; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_751 = 12'h2ef == csr_addr[11:0] ? reg_csr_751 : _GEN_750; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_752 = 12'h2f0 == csr_addr[11:0] ? reg_csr_752 : _GEN_751; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_753 = 12'h2f1 == csr_addr[11:0] ? reg_csr_753 : _GEN_752; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_754 = 12'h2f2 == csr_addr[11:0] ? reg_csr_754 : _GEN_753; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_755 = 12'h2f3 == csr_addr[11:0] ? reg_csr_755 : _GEN_754; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_756 = 12'h2f4 == csr_addr[11:0] ? reg_csr_756 : _GEN_755; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_757 = 12'h2f5 == csr_addr[11:0] ? reg_csr_757 : _GEN_756; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_758 = 12'h2f6 == csr_addr[11:0] ? reg_csr_758 : _GEN_757; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_759 = 12'h2f7 == csr_addr[11:0] ? reg_csr_759 : _GEN_758; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_760 = 12'h2f8 == csr_addr[11:0] ? reg_csr_760 : _GEN_759; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_761 = 12'h2f9 == csr_addr[11:0] ? reg_csr_761 : _GEN_760; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_762 = 12'h2fa == csr_addr[11:0] ? reg_csr_762 : _GEN_761; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_763 = 12'h2fb == csr_addr[11:0] ? reg_csr_763 : _GEN_762; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_764 = 12'h2fc == csr_addr[11:0] ? reg_csr_764 : _GEN_763; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_765 = 12'h2fd == csr_addr[11:0] ? reg_csr_765 : _GEN_764; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_766 = 12'h2fe == csr_addr[11:0] ? reg_csr_766 : _GEN_765; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_767 = 12'h2ff == csr_addr[11:0] ? reg_csr_767 : _GEN_766; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_768 = 12'h300 == csr_addr[11:0] ? reg_csr_768 : _GEN_767; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_769 = 12'h301 == csr_addr[11:0] ? reg_csr_769 : _GEN_768; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_770 = 12'h302 == csr_addr[11:0] ? reg_csr_770 : _GEN_769; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_771 = 12'h303 == csr_addr[11:0] ? reg_csr_771 : _GEN_770; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_772 = 12'h304 == csr_addr[11:0] ? reg_csr_772 : _GEN_771; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_773 = 12'h305 == csr_addr[11:0] ? reg_csr_773 : _GEN_772; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_774 = 12'h306 == csr_addr[11:0] ? reg_csr_774 : _GEN_773; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_775 = 12'h307 == csr_addr[11:0] ? reg_csr_775 : _GEN_774; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_776 = 12'h308 == csr_addr[11:0] ? reg_csr_776 : _GEN_775; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_777 = 12'h309 == csr_addr[11:0] ? reg_csr_777 : _GEN_776; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_778 = 12'h30a == csr_addr[11:0] ? reg_csr_778 : _GEN_777; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_779 = 12'h30b == csr_addr[11:0] ? reg_csr_779 : _GEN_778; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_780 = 12'h30c == csr_addr[11:0] ? reg_csr_780 : _GEN_779; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_781 = 12'h30d == csr_addr[11:0] ? reg_csr_781 : _GEN_780; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_782 = 12'h30e == csr_addr[11:0] ? reg_csr_782 : _GEN_781; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_783 = 12'h30f == csr_addr[11:0] ? reg_csr_783 : _GEN_782; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_784 = 12'h310 == csr_addr[11:0] ? reg_csr_784 : _GEN_783; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_785 = 12'h311 == csr_addr[11:0] ? reg_csr_785 : _GEN_784; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_786 = 12'h312 == csr_addr[11:0] ? reg_csr_786 : _GEN_785; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_787 = 12'h313 == csr_addr[11:0] ? reg_csr_787 : _GEN_786; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_788 = 12'h314 == csr_addr[11:0] ? reg_csr_788 : _GEN_787; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_789 = 12'h315 == csr_addr[11:0] ? reg_csr_789 : _GEN_788; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_790 = 12'h316 == csr_addr[11:0] ? reg_csr_790 : _GEN_789; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_791 = 12'h317 == csr_addr[11:0] ? reg_csr_791 : _GEN_790; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_792 = 12'h318 == csr_addr[11:0] ? reg_csr_792 : _GEN_791; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_793 = 12'h319 == csr_addr[11:0] ? reg_csr_793 : _GEN_792; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_794 = 12'h31a == csr_addr[11:0] ? reg_csr_794 : _GEN_793; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_795 = 12'h31b == csr_addr[11:0] ? reg_csr_795 : _GEN_794; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_796 = 12'h31c == csr_addr[11:0] ? reg_csr_796 : _GEN_795; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_797 = 12'h31d == csr_addr[11:0] ? reg_csr_797 : _GEN_796; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_798 = 12'h31e == csr_addr[11:0] ? reg_csr_798 : _GEN_797; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_799 = 12'h31f == csr_addr[11:0] ? reg_csr_799 : _GEN_798; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_800 = 12'h320 == csr_addr[11:0] ? reg_csr_800 : _GEN_799; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_801 = 12'h321 == csr_addr[11:0] ? reg_csr_801 : _GEN_800; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_802 = 12'h322 == csr_addr[11:0] ? reg_csr_802 : _GEN_801; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_803 = 12'h323 == csr_addr[11:0] ? reg_csr_803 : _GEN_802; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_804 = 12'h324 == csr_addr[11:0] ? reg_csr_804 : _GEN_803; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_805 = 12'h325 == csr_addr[11:0] ? reg_csr_805 : _GEN_804; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_806 = 12'h326 == csr_addr[11:0] ? reg_csr_806 : _GEN_805; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_807 = 12'h327 == csr_addr[11:0] ? reg_csr_807 : _GEN_806; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_808 = 12'h328 == csr_addr[11:0] ? reg_csr_808 : _GEN_807; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_809 = 12'h329 == csr_addr[11:0] ? reg_csr_809 : _GEN_808; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_810 = 12'h32a == csr_addr[11:0] ? reg_csr_810 : _GEN_809; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_811 = 12'h32b == csr_addr[11:0] ? reg_csr_811 : _GEN_810; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_812 = 12'h32c == csr_addr[11:0] ? reg_csr_812 : _GEN_811; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_813 = 12'h32d == csr_addr[11:0] ? reg_csr_813 : _GEN_812; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_814 = 12'h32e == csr_addr[11:0] ? reg_csr_814 : _GEN_813; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_815 = 12'h32f == csr_addr[11:0] ? reg_csr_815 : _GEN_814; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_816 = 12'h330 == csr_addr[11:0] ? reg_csr_816 : _GEN_815; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_817 = 12'h331 == csr_addr[11:0] ? reg_csr_817 : _GEN_816; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_818 = 12'h332 == csr_addr[11:0] ? reg_csr_818 : _GEN_817; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_819 = 12'h333 == csr_addr[11:0] ? reg_csr_819 : _GEN_818; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_820 = 12'h334 == csr_addr[11:0] ? reg_csr_820 : _GEN_819; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_821 = 12'h335 == csr_addr[11:0] ? reg_csr_821 : _GEN_820; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_822 = 12'h336 == csr_addr[11:0] ? reg_csr_822 : _GEN_821; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_823 = 12'h337 == csr_addr[11:0] ? reg_csr_823 : _GEN_822; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_824 = 12'h338 == csr_addr[11:0] ? reg_csr_824 : _GEN_823; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_825 = 12'h339 == csr_addr[11:0] ? reg_csr_825 : _GEN_824; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_826 = 12'h33a == csr_addr[11:0] ? reg_csr_826 : _GEN_825; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_827 = 12'h33b == csr_addr[11:0] ? reg_csr_827 : _GEN_826; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_828 = 12'h33c == csr_addr[11:0] ? reg_csr_828 : _GEN_827; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_829 = 12'h33d == csr_addr[11:0] ? reg_csr_829 : _GEN_828; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_830 = 12'h33e == csr_addr[11:0] ? reg_csr_830 : _GEN_829; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_831 = 12'h33f == csr_addr[11:0] ? reg_csr_831 : _GEN_830; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_832 = 12'h340 == csr_addr[11:0] ? reg_csr_832 : _GEN_831; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_833 = 12'h341 == csr_addr[11:0] ? reg_csr_833 : _GEN_832; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_834 = 12'h342 == csr_addr[11:0] ? reg_csr_834 : _GEN_833; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_835 = 12'h343 == csr_addr[11:0] ? reg_csr_835 : _GEN_834; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_836 = 12'h344 == csr_addr[11:0] ? reg_csr_836 : _GEN_835; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_837 = 12'h345 == csr_addr[11:0] ? reg_csr_837 : _GEN_836; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_838 = 12'h346 == csr_addr[11:0] ? reg_csr_838 : _GEN_837; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_839 = 12'h347 == csr_addr[11:0] ? reg_csr_839 : _GEN_838; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_840 = 12'h348 == csr_addr[11:0] ? reg_csr_840 : _GEN_839; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_841 = 12'h349 == csr_addr[11:0] ? reg_csr_841 : _GEN_840; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_842 = 12'h34a == csr_addr[11:0] ? reg_csr_842 : _GEN_841; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_843 = 12'h34b == csr_addr[11:0] ? reg_csr_843 : _GEN_842; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_844 = 12'h34c == csr_addr[11:0] ? reg_csr_844 : _GEN_843; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_845 = 12'h34d == csr_addr[11:0] ? reg_csr_845 : _GEN_844; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_846 = 12'h34e == csr_addr[11:0] ? reg_csr_846 : _GEN_845; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_847 = 12'h34f == csr_addr[11:0] ? reg_csr_847 : _GEN_846; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_848 = 12'h350 == csr_addr[11:0] ? reg_csr_848 : _GEN_847; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_849 = 12'h351 == csr_addr[11:0] ? reg_csr_849 : _GEN_848; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_850 = 12'h352 == csr_addr[11:0] ? reg_csr_850 : _GEN_849; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_851 = 12'h353 == csr_addr[11:0] ? reg_csr_851 : _GEN_850; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_852 = 12'h354 == csr_addr[11:0] ? reg_csr_852 : _GEN_851; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_853 = 12'h355 == csr_addr[11:0] ? reg_csr_853 : _GEN_852; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_854 = 12'h356 == csr_addr[11:0] ? reg_csr_854 : _GEN_853; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_855 = 12'h357 == csr_addr[11:0] ? reg_csr_855 : _GEN_854; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_856 = 12'h358 == csr_addr[11:0] ? reg_csr_856 : _GEN_855; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_857 = 12'h359 == csr_addr[11:0] ? reg_csr_857 : _GEN_856; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_858 = 12'h35a == csr_addr[11:0] ? reg_csr_858 : _GEN_857; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_859 = 12'h35b == csr_addr[11:0] ? reg_csr_859 : _GEN_858; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_860 = 12'h35c == csr_addr[11:0] ? reg_csr_860 : _GEN_859; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_861 = 12'h35d == csr_addr[11:0] ? reg_csr_861 : _GEN_860; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_862 = 12'h35e == csr_addr[11:0] ? reg_csr_862 : _GEN_861; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_863 = 12'h35f == csr_addr[11:0] ? reg_csr_863 : _GEN_862; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_864 = 12'h360 == csr_addr[11:0] ? reg_csr_864 : _GEN_863; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_865 = 12'h361 == csr_addr[11:0] ? reg_csr_865 : _GEN_864; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_866 = 12'h362 == csr_addr[11:0] ? reg_csr_866 : _GEN_865; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_867 = 12'h363 == csr_addr[11:0] ? reg_csr_867 : _GEN_866; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_868 = 12'h364 == csr_addr[11:0] ? reg_csr_868 : _GEN_867; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_869 = 12'h365 == csr_addr[11:0] ? reg_csr_869 : _GEN_868; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_870 = 12'h366 == csr_addr[11:0] ? reg_csr_870 : _GEN_869; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_871 = 12'h367 == csr_addr[11:0] ? reg_csr_871 : _GEN_870; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_872 = 12'h368 == csr_addr[11:0] ? reg_csr_872 : _GEN_871; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_873 = 12'h369 == csr_addr[11:0] ? reg_csr_873 : _GEN_872; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_874 = 12'h36a == csr_addr[11:0] ? reg_csr_874 : _GEN_873; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_875 = 12'h36b == csr_addr[11:0] ? reg_csr_875 : _GEN_874; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_876 = 12'h36c == csr_addr[11:0] ? reg_csr_876 : _GEN_875; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_877 = 12'h36d == csr_addr[11:0] ? reg_csr_877 : _GEN_876; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_878 = 12'h36e == csr_addr[11:0] ? reg_csr_878 : _GEN_877; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_879 = 12'h36f == csr_addr[11:0] ? reg_csr_879 : _GEN_878; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_880 = 12'h370 == csr_addr[11:0] ? reg_csr_880 : _GEN_879; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_881 = 12'h371 == csr_addr[11:0] ? reg_csr_881 : _GEN_880; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_882 = 12'h372 == csr_addr[11:0] ? reg_csr_882 : _GEN_881; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_883 = 12'h373 == csr_addr[11:0] ? reg_csr_883 : _GEN_882; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_884 = 12'h374 == csr_addr[11:0] ? reg_csr_884 : _GEN_883; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_885 = 12'h375 == csr_addr[11:0] ? reg_csr_885 : _GEN_884; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_886 = 12'h376 == csr_addr[11:0] ? reg_csr_886 : _GEN_885; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_887 = 12'h377 == csr_addr[11:0] ? reg_csr_887 : _GEN_886; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_888 = 12'h378 == csr_addr[11:0] ? reg_csr_888 : _GEN_887; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_889 = 12'h379 == csr_addr[11:0] ? reg_csr_889 : _GEN_888; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_890 = 12'h37a == csr_addr[11:0] ? reg_csr_890 : _GEN_889; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_891 = 12'h37b == csr_addr[11:0] ? reg_csr_891 : _GEN_890; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_892 = 12'h37c == csr_addr[11:0] ? reg_csr_892 : _GEN_891; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_893 = 12'h37d == csr_addr[11:0] ? reg_csr_893 : _GEN_892; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_894 = 12'h37e == csr_addr[11:0] ? reg_csr_894 : _GEN_893; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_895 = 12'h37f == csr_addr[11:0] ? reg_csr_895 : _GEN_894; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_896 = 12'h380 == csr_addr[11:0] ? reg_csr_896 : _GEN_895; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_897 = 12'h381 == csr_addr[11:0] ? reg_csr_897 : _GEN_896; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_898 = 12'h382 == csr_addr[11:0] ? reg_csr_898 : _GEN_897; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_899 = 12'h383 == csr_addr[11:0] ? reg_csr_899 : _GEN_898; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_900 = 12'h384 == csr_addr[11:0] ? reg_csr_900 : _GEN_899; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_901 = 12'h385 == csr_addr[11:0] ? reg_csr_901 : _GEN_900; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_902 = 12'h386 == csr_addr[11:0] ? reg_csr_902 : _GEN_901; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_903 = 12'h387 == csr_addr[11:0] ? reg_csr_903 : _GEN_902; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_904 = 12'h388 == csr_addr[11:0] ? reg_csr_904 : _GEN_903; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_905 = 12'h389 == csr_addr[11:0] ? reg_csr_905 : _GEN_904; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_906 = 12'h38a == csr_addr[11:0] ? reg_csr_906 : _GEN_905; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_907 = 12'h38b == csr_addr[11:0] ? reg_csr_907 : _GEN_906; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_908 = 12'h38c == csr_addr[11:0] ? reg_csr_908 : _GEN_907; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_909 = 12'h38d == csr_addr[11:0] ? reg_csr_909 : _GEN_908; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_910 = 12'h38e == csr_addr[11:0] ? reg_csr_910 : _GEN_909; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_911 = 12'h38f == csr_addr[11:0] ? reg_csr_911 : _GEN_910; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_912 = 12'h390 == csr_addr[11:0] ? reg_csr_912 : _GEN_911; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_913 = 12'h391 == csr_addr[11:0] ? reg_csr_913 : _GEN_912; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_914 = 12'h392 == csr_addr[11:0] ? reg_csr_914 : _GEN_913; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_915 = 12'h393 == csr_addr[11:0] ? reg_csr_915 : _GEN_914; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_916 = 12'h394 == csr_addr[11:0] ? reg_csr_916 : _GEN_915; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_917 = 12'h395 == csr_addr[11:0] ? reg_csr_917 : _GEN_916; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_918 = 12'h396 == csr_addr[11:0] ? reg_csr_918 : _GEN_917; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_919 = 12'h397 == csr_addr[11:0] ? reg_csr_919 : _GEN_918; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_920 = 12'h398 == csr_addr[11:0] ? reg_csr_920 : _GEN_919; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_921 = 12'h399 == csr_addr[11:0] ? reg_csr_921 : _GEN_920; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_922 = 12'h39a == csr_addr[11:0] ? reg_csr_922 : _GEN_921; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_923 = 12'h39b == csr_addr[11:0] ? reg_csr_923 : _GEN_922; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_924 = 12'h39c == csr_addr[11:0] ? reg_csr_924 : _GEN_923; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_925 = 12'h39d == csr_addr[11:0] ? reg_csr_925 : _GEN_924; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_926 = 12'h39e == csr_addr[11:0] ? reg_csr_926 : _GEN_925; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_927 = 12'h39f == csr_addr[11:0] ? reg_csr_927 : _GEN_926; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_928 = 12'h3a0 == csr_addr[11:0] ? reg_csr_928 : _GEN_927; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_929 = 12'h3a1 == csr_addr[11:0] ? reg_csr_929 : _GEN_928; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_930 = 12'h3a2 == csr_addr[11:0] ? reg_csr_930 : _GEN_929; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_931 = 12'h3a3 == csr_addr[11:0] ? reg_csr_931 : _GEN_930; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_932 = 12'h3a4 == csr_addr[11:0] ? reg_csr_932 : _GEN_931; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_933 = 12'h3a5 == csr_addr[11:0] ? reg_csr_933 : _GEN_932; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_934 = 12'h3a6 == csr_addr[11:0] ? reg_csr_934 : _GEN_933; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_935 = 12'h3a7 == csr_addr[11:0] ? reg_csr_935 : _GEN_934; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_936 = 12'h3a8 == csr_addr[11:0] ? reg_csr_936 : _GEN_935; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_937 = 12'h3a9 == csr_addr[11:0] ? reg_csr_937 : _GEN_936; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_938 = 12'h3aa == csr_addr[11:0] ? reg_csr_938 : _GEN_937; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_939 = 12'h3ab == csr_addr[11:0] ? reg_csr_939 : _GEN_938; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_940 = 12'h3ac == csr_addr[11:0] ? reg_csr_940 : _GEN_939; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_941 = 12'h3ad == csr_addr[11:0] ? reg_csr_941 : _GEN_940; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_942 = 12'h3ae == csr_addr[11:0] ? reg_csr_942 : _GEN_941; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_943 = 12'h3af == csr_addr[11:0] ? reg_csr_943 : _GEN_942; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_944 = 12'h3b0 == csr_addr[11:0] ? reg_csr_944 : _GEN_943; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_945 = 12'h3b1 == csr_addr[11:0] ? reg_csr_945 : _GEN_944; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_946 = 12'h3b2 == csr_addr[11:0] ? reg_csr_946 : _GEN_945; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_947 = 12'h3b3 == csr_addr[11:0] ? reg_csr_947 : _GEN_946; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_948 = 12'h3b4 == csr_addr[11:0] ? reg_csr_948 : _GEN_947; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_949 = 12'h3b5 == csr_addr[11:0] ? reg_csr_949 : _GEN_948; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_950 = 12'h3b6 == csr_addr[11:0] ? reg_csr_950 : _GEN_949; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_951 = 12'h3b7 == csr_addr[11:0] ? reg_csr_951 : _GEN_950; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_952 = 12'h3b8 == csr_addr[11:0] ? reg_csr_952 : _GEN_951; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_953 = 12'h3b9 == csr_addr[11:0] ? reg_csr_953 : _GEN_952; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_954 = 12'h3ba == csr_addr[11:0] ? reg_csr_954 : _GEN_953; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_955 = 12'h3bb == csr_addr[11:0] ? reg_csr_955 : _GEN_954; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_956 = 12'h3bc == csr_addr[11:0] ? reg_csr_956 : _GEN_955; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_957 = 12'h3bd == csr_addr[11:0] ? reg_csr_957 : _GEN_956; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_958 = 12'h3be == csr_addr[11:0] ? reg_csr_958 : _GEN_957; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_959 = 12'h3bf == csr_addr[11:0] ? reg_csr_959 : _GEN_958; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_960 = 12'h3c0 == csr_addr[11:0] ? reg_csr_960 : _GEN_959; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_961 = 12'h3c1 == csr_addr[11:0] ? reg_csr_961 : _GEN_960; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_962 = 12'h3c2 == csr_addr[11:0] ? reg_csr_962 : _GEN_961; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_963 = 12'h3c3 == csr_addr[11:0] ? reg_csr_963 : _GEN_962; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_964 = 12'h3c4 == csr_addr[11:0] ? reg_csr_964 : _GEN_963; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_965 = 12'h3c5 == csr_addr[11:0] ? reg_csr_965 : _GEN_964; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_966 = 12'h3c6 == csr_addr[11:0] ? reg_csr_966 : _GEN_965; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_967 = 12'h3c7 == csr_addr[11:0] ? reg_csr_967 : _GEN_966; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_968 = 12'h3c8 == csr_addr[11:0] ? reg_csr_968 : _GEN_967; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_969 = 12'h3c9 == csr_addr[11:0] ? reg_csr_969 : _GEN_968; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_970 = 12'h3ca == csr_addr[11:0] ? reg_csr_970 : _GEN_969; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_971 = 12'h3cb == csr_addr[11:0] ? reg_csr_971 : _GEN_970; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_972 = 12'h3cc == csr_addr[11:0] ? reg_csr_972 : _GEN_971; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_973 = 12'h3cd == csr_addr[11:0] ? reg_csr_973 : _GEN_972; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_974 = 12'h3ce == csr_addr[11:0] ? reg_csr_974 : _GEN_973; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_975 = 12'h3cf == csr_addr[11:0] ? reg_csr_975 : _GEN_974; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_976 = 12'h3d0 == csr_addr[11:0] ? reg_csr_976 : _GEN_975; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_977 = 12'h3d1 == csr_addr[11:0] ? reg_csr_977 : _GEN_976; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_978 = 12'h3d2 == csr_addr[11:0] ? reg_csr_978 : _GEN_977; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_979 = 12'h3d3 == csr_addr[11:0] ? reg_csr_979 : _GEN_978; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_980 = 12'h3d4 == csr_addr[11:0] ? reg_csr_980 : _GEN_979; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_981 = 12'h3d5 == csr_addr[11:0] ? reg_csr_981 : _GEN_980; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_982 = 12'h3d6 == csr_addr[11:0] ? reg_csr_982 : _GEN_981; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_983 = 12'h3d7 == csr_addr[11:0] ? reg_csr_983 : _GEN_982; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_984 = 12'h3d8 == csr_addr[11:0] ? reg_csr_984 : _GEN_983; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_985 = 12'h3d9 == csr_addr[11:0] ? reg_csr_985 : _GEN_984; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_986 = 12'h3da == csr_addr[11:0] ? reg_csr_986 : _GEN_985; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_987 = 12'h3db == csr_addr[11:0] ? reg_csr_987 : _GEN_986; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_988 = 12'h3dc == csr_addr[11:0] ? reg_csr_988 : _GEN_987; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_989 = 12'h3dd == csr_addr[11:0] ? reg_csr_989 : _GEN_988; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_990 = 12'h3de == csr_addr[11:0] ? reg_csr_990 : _GEN_989; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_991 = 12'h3df == csr_addr[11:0] ? reg_csr_991 : _GEN_990; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_992 = 12'h3e0 == csr_addr[11:0] ? reg_csr_992 : _GEN_991; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_993 = 12'h3e1 == csr_addr[11:0] ? reg_csr_993 : _GEN_992; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_994 = 12'h3e2 == csr_addr[11:0] ? reg_csr_994 : _GEN_993; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_995 = 12'h3e3 == csr_addr[11:0] ? reg_csr_995 : _GEN_994; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_996 = 12'h3e4 == csr_addr[11:0] ? reg_csr_996 : _GEN_995; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_997 = 12'h3e5 == csr_addr[11:0] ? reg_csr_997 : _GEN_996; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_998 = 12'h3e6 == csr_addr[11:0] ? reg_csr_998 : _GEN_997; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_999 = 12'h3e7 == csr_addr[11:0] ? reg_csr_999 : _GEN_998; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1000 = 12'h3e8 == csr_addr[11:0] ? reg_csr_1000 : _GEN_999; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1001 = 12'h3e9 == csr_addr[11:0] ? reg_csr_1001 : _GEN_1000; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1002 = 12'h3ea == csr_addr[11:0] ? reg_csr_1002 : _GEN_1001; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1003 = 12'h3eb == csr_addr[11:0] ? reg_csr_1003 : _GEN_1002; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1004 = 12'h3ec == csr_addr[11:0] ? reg_csr_1004 : _GEN_1003; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1005 = 12'h3ed == csr_addr[11:0] ? reg_csr_1005 : _GEN_1004; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1006 = 12'h3ee == csr_addr[11:0] ? reg_csr_1006 : _GEN_1005; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1007 = 12'h3ef == csr_addr[11:0] ? reg_csr_1007 : _GEN_1006; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1008 = 12'h3f0 == csr_addr[11:0] ? reg_csr_1008 : _GEN_1007; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1009 = 12'h3f1 == csr_addr[11:0] ? reg_csr_1009 : _GEN_1008; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1010 = 12'h3f2 == csr_addr[11:0] ? reg_csr_1010 : _GEN_1009; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1011 = 12'h3f3 == csr_addr[11:0] ? reg_csr_1011 : _GEN_1010; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1012 = 12'h3f4 == csr_addr[11:0] ? reg_csr_1012 : _GEN_1011; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1013 = 12'h3f5 == csr_addr[11:0] ? reg_csr_1013 : _GEN_1012; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1014 = 12'h3f6 == csr_addr[11:0] ? reg_csr_1014 : _GEN_1013; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1015 = 12'h3f7 == csr_addr[11:0] ? reg_csr_1015 : _GEN_1014; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1016 = 12'h3f8 == csr_addr[11:0] ? reg_csr_1016 : _GEN_1015; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1017 = 12'h3f9 == csr_addr[11:0] ? reg_csr_1017 : _GEN_1016; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1018 = 12'h3fa == csr_addr[11:0] ? reg_csr_1018 : _GEN_1017; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1019 = 12'h3fb == csr_addr[11:0] ? reg_csr_1019 : _GEN_1018; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1020 = 12'h3fc == csr_addr[11:0] ? reg_csr_1020 : _GEN_1019; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1021 = 12'h3fd == csr_addr[11:0] ? reg_csr_1021 : _GEN_1020; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1022 = 12'h3fe == csr_addr[11:0] ? reg_csr_1022 : _GEN_1021; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1023 = 12'h3ff == csr_addr[11:0] ? reg_csr_1023 : _GEN_1022; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1024 = 12'h400 == csr_addr[11:0] ? reg_csr_1024 : _GEN_1023; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1025 = 12'h401 == csr_addr[11:0] ? reg_csr_1025 : _GEN_1024; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1026 = 12'h402 == csr_addr[11:0] ? reg_csr_1026 : _GEN_1025; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1027 = 12'h403 == csr_addr[11:0] ? reg_csr_1027 : _GEN_1026; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1028 = 12'h404 == csr_addr[11:0] ? reg_csr_1028 : _GEN_1027; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1029 = 12'h405 == csr_addr[11:0] ? reg_csr_1029 : _GEN_1028; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1030 = 12'h406 == csr_addr[11:0] ? reg_csr_1030 : _GEN_1029; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1031 = 12'h407 == csr_addr[11:0] ? reg_csr_1031 : _GEN_1030; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1032 = 12'h408 == csr_addr[11:0] ? reg_csr_1032 : _GEN_1031; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1033 = 12'h409 == csr_addr[11:0] ? reg_csr_1033 : _GEN_1032; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1034 = 12'h40a == csr_addr[11:0] ? reg_csr_1034 : _GEN_1033; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1035 = 12'h40b == csr_addr[11:0] ? reg_csr_1035 : _GEN_1034; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1036 = 12'h40c == csr_addr[11:0] ? reg_csr_1036 : _GEN_1035; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1037 = 12'h40d == csr_addr[11:0] ? reg_csr_1037 : _GEN_1036; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1038 = 12'h40e == csr_addr[11:0] ? reg_csr_1038 : _GEN_1037; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1039 = 12'h40f == csr_addr[11:0] ? reg_csr_1039 : _GEN_1038; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1040 = 12'h410 == csr_addr[11:0] ? reg_csr_1040 : _GEN_1039; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1041 = 12'h411 == csr_addr[11:0] ? reg_csr_1041 : _GEN_1040; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1042 = 12'h412 == csr_addr[11:0] ? reg_csr_1042 : _GEN_1041; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1043 = 12'h413 == csr_addr[11:0] ? reg_csr_1043 : _GEN_1042; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1044 = 12'h414 == csr_addr[11:0] ? reg_csr_1044 : _GEN_1043; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1045 = 12'h415 == csr_addr[11:0] ? reg_csr_1045 : _GEN_1044; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1046 = 12'h416 == csr_addr[11:0] ? reg_csr_1046 : _GEN_1045; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1047 = 12'h417 == csr_addr[11:0] ? reg_csr_1047 : _GEN_1046; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1048 = 12'h418 == csr_addr[11:0] ? reg_csr_1048 : _GEN_1047; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1049 = 12'h419 == csr_addr[11:0] ? reg_csr_1049 : _GEN_1048; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1050 = 12'h41a == csr_addr[11:0] ? reg_csr_1050 : _GEN_1049; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1051 = 12'h41b == csr_addr[11:0] ? reg_csr_1051 : _GEN_1050; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1052 = 12'h41c == csr_addr[11:0] ? reg_csr_1052 : _GEN_1051; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1053 = 12'h41d == csr_addr[11:0] ? reg_csr_1053 : _GEN_1052; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1054 = 12'h41e == csr_addr[11:0] ? reg_csr_1054 : _GEN_1053; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1055 = 12'h41f == csr_addr[11:0] ? reg_csr_1055 : _GEN_1054; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1056 = 12'h420 == csr_addr[11:0] ? reg_csr_1056 : _GEN_1055; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1057 = 12'h421 == csr_addr[11:0] ? reg_csr_1057 : _GEN_1056; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1058 = 12'h422 == csr_addr[11:0] ? reg_csr_1058 : _GEN_1057; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1059 = 12'h423 == csr_addr[11:0] ? reg_csr_1059 : _GEN_1058; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1060 = 12'h424 == csr_addr[11:0] ? reg_csr_1060 : _GEN_1059; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1061 = 12'h425 == csr_addr[11:0] ? reg_csr_1061 : _GEN_1060; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1062 = 12'h426 == csr_addr[11:0] ? reg_csr_1062 : _GEN_1061; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1063 = 12'h427 == csr_addr[11:0] ? reg_csr_1063 : _GEN_1062; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1064 = 12'h428 == csr_addr[11:0] ? reg_csr_1064 : _GEN_1063; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1065 = 12'h429 == csr_addr[11:0] ? reg_csr_1065 : _GEN_1064; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1066 = 12'h42a == csr_addr[11:0] ? reg_csr_1066 : _GEN_1065; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1067 = 12'h42b == csr_addr[11:0] ? reg_csr_1067 : _GEN_1066; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1068 = 12'h42c == csr_addr[11:0] ? reg_csr_1068 : _GEN_1067; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1069 = 12'h42d == csr_addr[11:0] ? reg_csr_1069 : _GEN_1068; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1070 = 12'h42e == csr_addr[11:0] ? reg_csr_1070 : _GEN_1069; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1071 = 12'h42f == csr_addr[11:0] ? reg_csr_1071 : _GEN_1070; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1072 = 12'h430 == csr_addr[11:0] ? reg_csr_1072 : _GEN_1071; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1073 = 12'h431 == csr_addr[11:0] ? reg_csr_1073 : _GEN_1072; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1074 = 12'h432 == csr_addr[11:0] ? reg_csr_1074 : _GEN_1073; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1075 = 12'h433 == csr_addr[11:0] ? reg_csr_1075 : _GEN_1074; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1076 = 12'h434 == csr_addr[11:0] ? reg_csr_1076 : _GEN_1075; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1077 = 12'h435 == csr_addr[11:0] ? reg_csr_1077 : _GEN_1076; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1078 = 12'h436 == csr_addr[11:0] ? reg_csr_1078 : _GEN_1077; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1079 = 12'h437 == csr_addr[11:0] ? reg_csr_1079 : _GEN_1078; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1080 = 12'h438 == csr_addr[11:0] ? reg_csr_1080 : _GEN_1079; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1081 = 12'h439 == csr_addr[11:0] ? reg_csr_1081 : _GEN_1080; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1082 = 12'h43a == csr_addr[11:0] ? reg_csr_1082 : _GEN_1081; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1083 = 12'h43b == csr_addr[11:0] ? reg_csr_1083 : _GEN_1082; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1084 = 12'h43c == csr_addr[11:0] ? reg_csr_1084 : _GEN_1083; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1085 = 12'h43d == csr_addr[11:0] ? reg_csr_1085 : _GEN_1084; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1086 = 12'h43e == csr_addr[11:0] ? reg_csr_1086 : _GEN_1085; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1087 = 12'h43f == csr_addr[11:0] ? reg_csr_1087 : _GEN_1086; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1088 = 12'h440 == csr_addr[11:0] ? reg_csr_1088 : _GEN_1087; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1089 = 12'h441 == csr_addr[11:0] ? reg_csr_1089 : _GEN_1088; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1090 = 12'h442 == csr_addr[11:0] ? reg_csr_1090 : _GEN_1089; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1091 = 12'h443 == csr_addr[11:0] ? reg_csr_1091 : _GEN_1090; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1092 = 12'h444 == csr_addr[11:0] ? reg_csr_1092 : _GEN_1091; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1093 = 12'h445 == csr_addr[11:0] ? reg_csr_1093 : _GEN_1092; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1094 = 12'h446 == csr_addr[11:0] ? reg_csr_1094 : _GEN_1093; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1095 = 12'h447 == csr_addr[11:0] ? reg_csr_1095 : _GEN_1094; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1096 = 12'h448 == csr_addr[11:0] ? reg_csr_1096 : _GEN_1095; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1097 = 12'h449 == csr_addr[11:0] ? reg_csr_1097 : _GEN_1096; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1098 = 12'h44a == csr_addr[11:0] ? reg_csr_1098 : _GEN_1097; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1099 = 12'h44b == csr_addr[11:0] ? reg_csr_1099 : _GEN_1098; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1100 = 12'h44c == csr_addr[11:0] ? reg_csr_1100 : _GEN_1099; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1101 = 12'h44d == csr_addr[11:0] ? reg_csr_1101 : _GEN_1100; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1102 = 12'h44e == csr_addr[11:0] ? reg_csr_1102 : _GEN_1101; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1103 = 12'h44f == csr_addr[11:0] ? reg_csr_1103 : _GEN_1102; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1104 = 12'h450 == csr_addr[11:0] ? reg_csr_1104 : _GEN_1103; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1105 = 12'h451 == csr_addr[11:0] ? reg_csr_1105 : _GEN_1104; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1106 = 12'h452 == csr_addr[11:0] ? reg_csr_1106 : _GEN_1105; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1107 = 12'h453 == csr_addr[11:0] ? reg_csr_1107 : _GEN_1106; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1108 = 12'h454 == csr_addr[11:0] ? reg_csr_1108 : _GEN_1107; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1109 = 12'h455 == csr_addr[11:0] ? reg_csr_1109 : _GEN_1108; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1110 = 12'h456 == csr_addr[11:0] ? reg_csr_1110 : _GEN_1109; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1111 = 12'h457 == csr_addr[11:0] ? reg_csr_1111 : _GEN_1110; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1112 = 12'h458 == csr_addr[11:0] ? reg_csr_1112 : _GEN_1111; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1113 = 12'h459 == csr_addr[11:0] ? reg_csr_1113 : _GEN_1112; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1114 = 12'h45a == csr_addr[11:0] ? reg_csr_1114 : _GEN_1113; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1115 = 12'h45b == csr_addr[11:0] ? reg_csr_1115 : _GEN_1114; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1116 = 12'h45c == csr_addr[11:0] ? reg_csr_1116 : _GEN_1115; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1117 = 12'h45d == csr_addr[11:0] ? reg_csr_1117 : _GEN_1116; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1118 = 12'h45e == csr_addr[11:0] ? reg_csr_1118 : _GEN_1117; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1119 = 12'h45f == csr_addr[11:0] ? reg_csr_1119 : _GEN_1118; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1120 = 12'h460 == csr_addr[11:0] ? reg_csr_1120 : _GEN_1119; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1121 = 12'h461 == csr_addr[11:0] ? reg_csr_1121 : _GEN_1120; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1122 = 12'h462 == csr_addr[11:0] ? reg_csr_1122 : _GEN_1121; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1123 = 12'h463 == csr_addr[11:0] ? reg_csr_1123 : _GEN_1122; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1124 = 12'h464 == csr_addr[11:0] ? reg_csr_1124 : _GEN_1123; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1125 = 12'h465 == csr_addr[11:0] ? reg_csr_1125 : _GEN_1124; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1126 = 12'h466 == csr_addr[11:0] ? reg_csr_1126 : _GEN_1125; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1127 = 12'h467 == csr_addr[11:0] ? reg_csr_1127 : _GEN_1126; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1128 = 12'h468 == csr_addr[11:0] ? reg_csr_1128 : _GEN_1127; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1129 = 12'h469 == csr_addr[11:0] ? reg_csr_1129 : _GEN_1128; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1130 = 12'h46a == csr_addr[11:0] ? reg_csr_1130 : _GEN_1129; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1131 = 12'h46b == csr_addr[11:0] ? reg_csr_1131 : _GEN_1130; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1132 = 12'h46c == csr_addr[11:0] ? reg_csr_1132 : _GEN_1131; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1133 = 12'h46d == csr_addr[11:0] ? reg_csr_1133 : _GEN_1132; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1134 = 12'h46e == csr_addr[11:0] ? reg_csr_1134 : _GEN_1133; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1135 = 12'h46f == csr_addr[11:0] ? reg_csr_1135 : _GEN_1134; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1136 = 12'h470 == csr_addr[11:0] ? reg_csr_1136 : _GEN_1135; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1137 = 12'h471 == csr_addr[11:0] ? reg_csr_1137 : _GEN_1136; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1138 = 12'h472 == csr_addr[11:0] ? reg_csr_1138 : _GEN_1137; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1139 = 12'h473 == csr_addr[11:0] ? reg_csr_1139 : _GEN_1138; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1140 = 12'h474 == csr_addr[11:0] ? reg_csr_1140 : _GEN_1139; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1141 = 12'h475 == csr_addr[11:0] ? reg_csr_1141 : _GEN_1140; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1142 = 12'h476 == csr_addr[11:0] ? reg_csr_1142 : _GEN_1141; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1143 = 12'h477 == csr_addr[11:0] ? reg_csr_1143 : _GEN_1142; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1144 = 12'h478 == csr_addr[11:0] ? reg_csr_1144 : _GEN_1143; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1145 = 12'h479 == csr_addr[11:0] ? reg_csr_1145 : _GEN_1144; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1146 = 12'h47a == csr_addr[11:0] ? reg_csr_1146 : _GEN_1145; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1147 = 12'h47b == csr_addr[11:0] ? reg_csr_1147 : _GEN_1146; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1148 = 12'h47c == csr_addr[11:0] ? reg_csr_1148 : _GEN_1147; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1149 = 12'h47d == csr_addr[11:0] ? reg_csr_1149 : _GEN_1148; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1150 = 12'h47e == csr_addr[11:0] ? reg_csr_1150 : _GEN_1149; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1151 = 12'h47f == csr_addr[11:0] ? reg_csr_1151 : _GEN_1150; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1152 = 12'h480 == csr_addr[11:0] ? reg_csr_1152 : _GEN_1151; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1153 = 12'h481 == csr_addr[11:0] ? reg_csr_1153 : _GEN_1152; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1154 = 12'h482 == csr_addr[11:0] ? reg_csr_1154 : _GEN_1153; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1155 = 12'h483 == csr_addr[11:0] ? reg_csr_1155 : _GEN_1154; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1156 = 12'h484 == csr_addr[11:0] ? reg_csr_1156 : _GEN_1155; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1157 = 12'h485 == csr_addr[11:0] ? reg_csr_1157 : _GEN_1156; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1158 = 12'h486 == csr_addr[11:0] ? reg_csr_1158 : _GEN_1157; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1159 = 12'h487 == csr_addr[11:0] ? reg_csr_1159 : _GEN_1158; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1160 = 12'h488 == csr_addr[11:0] ? reg_csr_1160 : _GEN_1159; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1161 = 12'h489 == csr_addr[11:0] ? reg_csr_1161 : _GEN_1160; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1162 = 12'h48a == csr_addr[11:0] ? reg_csr_1162 : _GEN_1161; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1163 = 12'h48b == csr_addr[11:0] ? reg_csr_1163 : _GEN_1162; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1164 = 12'h48c == csr_addr[11:0] ? reg_csr_1164 : _GEN_1163; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1165 = 12'h48d == csr_addr[11:0] ? reg_csr_1165 : _GEN_1164; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1166 = 12'h48e == csr_addr[11:0] ? reg_csr_1166 : _GEN_1165; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1167 = 12'h48f == csr_addr[11:0] ? reg_csr_1167 : _GEN_1166; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1168 = 12'h490 == csr_addr[11:0] ? reg_csr_1168 : _GEN_1167; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1169 = 12'h491 == csr_addr[11:0] ? reg_csr_1169 : _GEN_1168; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1170 = 12'h492 == csr_addr[11:0] ? reg_csr_1170 : _GEN_1169; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1171 = 12'h493 == csr_addr[11:0] ? reg_csr_1171 : _GEN_1170; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1172 = 12'h494 == csr_addr[11:0] ? reg_csr_1172 : _GEN_1171; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1173 = 12'h495 == csr_addr[11:0] ? reg_csr_1173 : _GEN_1172; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1174 = 12'h496 == csr_addr[11:0] ? reg_csr_1174 : _GEN_1173; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1175 = 12'h497 == csr_addr[11:0] ? reg_csr_1175 : _GEN_1174; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1176 = 12'h498 == csr_addr[11:0] ? reg_csr_1176 : _GEN_1175; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1177 = 12'h499 == csr_addr[11:0] ? reg_csr_1177 : _GEN_1176; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1178 = 12'h49a == csr_addr[11:0] ? reg_csr_1178 : _GEN_1177; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1179 = 12'h49b == csr_addr[11:0] ? reg_csr_1179 : _GEN_1178; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1180 = 12'h49c == csr_addr[11:0] ? reg_csr_1180 : _GEN_1179; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1181 = 12'h49d == csr_addr[11:0] ? reg_csr_1181 : _GEN_1180; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1182 = 12'h49e == csr_addr[11:0] ? reg_csr_1182 : _GEN_1181; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1183 = 12'h49f == csr_addr[11:0] ? reg_csr_1183 : _GEN_1182; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1184 = 12'h4a0 == csr_addr[11:0] ? reg_csr_1184 : _GEN_1183; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1185 = 12'h4a1 == csr_addr[11:0] ? reg_csr_1185 : _GEN_1184; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1186 = 12'h4a2 == csr_addr[11:0] ? reg_csr_1186 : _GEN_1185; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1187 = 12'h4a3 == csr_addr[11:0] ? reg_csr_1187 : _GEN_1186; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1188 = 12'h4a4 == csr_addr[11:0] ? reg_csr_1188 : _GEN_1187; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1189 = 12'h4a5 == csr_addr[11:0] ? reg_csr_1189 : _GEN_1188; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1190 = 12'h4a6 == csr_addr[11:0] ? reg_csr_1190 : _GEN_1189; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1191 = 12'h4a7 == csr_addr[11:0] ? reg_csr_1191 : _GEN_1190; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1192 = 12'h4a8 == csr_addr[11:0] ? reg_csr_1192 : _GEN_1191; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1193 = 12'h4a9 == csr_addr[11:0] ? reg_csr_1193 : _GEN_1192; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1194 = 12'h4aa == csr_addr[11:0] ? reg_csr_1194 : _GEN_1193; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1195 = 12'h4ab == csr_addr[11:0] ? reg_csr_1195 : _GEN_1194; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1196 = 12'h4ac == csr_addr[11:0] ? reg_csr_1196 : _GEN_1195; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1197 = 12'h4ad == csr_addr[11:0] ? reg_csr_1197 : _GEN_1196; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1198 = 12'h4ae == csr_addr[11:0] ? reg_csr_1198 : _GEN_1197; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1199 = 12'h4af == csr_addr[11:0] ? reg_csr_1199 : _GEN_1198; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1200 = 12'h4b0 == csr_addr[11:0] ? reg_csr_1200 : _GEN_1199; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1201 = 12'h4b1 == csr_addr[11:0] ? reg_csr_1201 : _GEN_1200; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1202 = 12'h4b2 == csr_addr[11:0] ? reg_csr_1202 : _GEN_1201; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1203 = 12'h4b3 == csr_addr[11:0] ? reg_csr_1203 : _GEN_1202; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1204 = 12'h4b4 == csr_addr[11:0] ? reg_csr_1204 : _GEN_1203; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1205 = 12'h4b5 == csr_addr[11:0] ? reg_csr_1205 : _GEN_1204; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1206 = 12'h4b6 == csr_addr[11:0] ? reg_csr_1206 : _GEN_1205; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1207 = 12'h4b7 == csr_addr[11:0] ? reg_csr_1207 : _GEN_1206; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1208 = 12'h4b8 == csr_addr[11:0] ? reg_csr_1208 : _GEN_1207; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1209 = 12'h4b9 == csr_addr[11:0] ? reg_csr_1209 : _GEN_1208; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1210 = 12'h4ba == csr_addr[11:0] ? reg_csr_1210 : _GEN_1209; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1211 = 12'h4bb == csr_addr[11:0] ? reg_csr_1211 : _GEN_1210; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1212 = 12'h4bc == csr_addr[11:0] ? reg_csr_1212 : _GEN_1211; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1213 = 12'h4bd == csr_addr[11:0] ? reg_csr_1213 : _GEN_1212; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1214 = 12'h4be == csr_addr[11:0] ? reg_csr_1214 : _GEN_1213; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1215 = 12'h4bf == csr_addr[11:0] ? reg_csr_1215 : _GEN_1214; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1216 = 12'h4c0 == csr_addr[11:0] ? reg_csr_1216 : _GEN_1215; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1217 = 12'h4c1 == csr_addr[11:0] ? reg_csr_1217 : _GEN_1216; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1218 = 12'h4c2 == csr_addr[11:0] ? reg_csr_1218 : _GEN_1217; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1219 = 12'h4c3 == csr_addr[11:0] ? reg_csr_1219 : _GEN_1218; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1220 = 12'h4c4 == csr_addr[11:0] ? reg_csr_1220 : _GEN_1219; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1221 = 12'h4c5 == csr_addr[11:0] ? reg_csr_1221 : _GEN_1220; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1222 = 12'h4c6 == csr_addr[11:0] ? reg_csr_1222 : _GEN_1221; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1223 = 12'h4c7 == csr_addr[11:0] ? reg_csr_1223 : _GEN_1222; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1224 = 12'h4c8 == csr_addr[11:0] ? reg_csr_1224 : _GEN_1223; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1225 = 12'h4c9 == csr_addr[11:0] ? reg_csr_1225 : _GEN_1224; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1226 = 12'h4ca == csr_addr[11:0] ? reg_csr_1226 : _GEN_1225; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1227 = 12'h4cb == csr_addr[11:0] ? reg_csr_1227 : _GEN_1226; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1228 = 12'h4cc == csr_addr[11:0] ? reg_csr_1228 : _GEN_1227; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1229 = 12'h4cd == csr_addr[11:0] ? reg_csr_1229 : _GEN_1228; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1230 = 12'h4ce == csr_addr[11:0] ? reg_csr_1230 : _GEN_1229; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1231 = 12'h4cf == csr_addr[11:0] ? reg_csr_1231 : _GEN_1230; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1232 = 12'h4d0 == csr_addr[11:0] ? reg_csr_1232 : _GEN_1231; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1233 = 12'h4d1 == csr_addr[11:0] ? reg_csr_1233 : _GEN_1232; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1234 = 12'h4d2 == csr_addr[11:0] ? reg_csr_1234 : _GEN_1233; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1235 = 12'h4d3 == csr_addr[11:0] ? reg_csr_1235 : _GEN_1234; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1236 = 12'h4d4 == csr_addr[11:0] ? reg_csr_1236 : _GEN_1235; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1237 = 12'h4d5 == csr_addr[11:0] ? reg_csr_1237 : _GEN_1236; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1238 = 12'h4d6 == csr_addr[11:0] ? reg_csr_1238 : _GEN_1237; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1239 = 12'h4d7 == csr_addr[11:0] ? reg_csr_1239 : _GEN_1238; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1240 = 12'h4d8 == csr_addr[11:0] ? reg_csr_1240 : _GEN_1239; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1241 = 12'h4d9 == csr_addr[11:0] ? reg_csr_1241 : _GEN_1240; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1242 = 12'h4da == csr_addr[11:0] ? reg_csr_1242 : _GEN_1241; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1243 = 12'h4db == csr_addr[11:0] ? reg_csr_1243 : _GEN_1242; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1244 = 12'h4dc == csr_addr[11:0] ? reg_csr_1244 : _GEN_1243; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1245 = 12'h4dd == csr_addr[11:0] ? reg_csr_1245 : _GEN_1244; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1246 = 12'h4de == csr_addr[11:0] ? reg_csr_1246 : _GEN_1245; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1247 = 12'h4df == csr_addr[11:0] ? reg_csr_1247 : _GEN_1246; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1248 = 12'h4e0 == csr_addr[11:0] ? reg_csr_1248 : _GEN_1247; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1249 = 12'h4e1 == csr_addr[11:0] ? reg_csr_1249 : _GEN_1248; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1250 = 12'h4e2 == csr_addr[11:0] ? reg_csr_1250 : _GEN_1249; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1251 = 12'h4e3 == csr_addr[11:0] ? reg_csr_1251 : _GEN_1250; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1252 = 12'h4e4 == csr_addr[11:0] ? reg_csr_1252 : _GEN_1251; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1253 = 12'h4e5 == csr_addr[11:0] ? reg_csr_1253 : _GEN_1252; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1254 = 12'h4e6 == csr_addr[11:0] ? reg_csr_1254 : _GEN_1253; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1255 = 12'h4e7 == csr_addr[11:0] ? reg_csr_1255 : _GEN_1254; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1256 = 12'h4e8 == csr_addr[11:0] ? reg_csr_1256 : _GEN_1255; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1257 = 12'h4e9 == csr_addr[11:0] ? reg_csr_1257 : _GEN_1256; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1258 = 12'h4ea == csr_addr[11:0] ? reg_csr_1258 : _GEN_1257; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1259 = 12'h4eb == csr_addr[11:0] ? reg_csr_1259 : _GEN_1258; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1260 = 12'h4ec == csr_addr[11:0] ? reg_csr_1260 : _GEN_1259; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1261 = 12'h4ed == csr_addr[11:0] ? reg_csr_1261 : _GEN_1260; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1262 = 12'h4ee == csr_addr[11:0] ? reg_csr_1262 : _GEN_1261; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1263 = 12'h4ef == csr_addr[11:0] ? reg_csr_1263 : _GEN_1262; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1264 = 12'h4f0 == csr_addr[11:0] ? reg_csr_1264 : _GEN_1263; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1265 = 12'h4f1 == csr_addr[11:0] ? reg_csr_1265 : _GEN_1264; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1266 = 12'h4f2 == csr_addr[11:0] ? reg_csr_1266 : _GEN_1265; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1267 = 12'h4f3 == csr_addr[11:0] ? reg_csr_1267 : _GEN_1266; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1268 = 12'h4f4 == csr_addr[11:0] ? reg_csr_1268 : _GEN_1267; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1269 = 12'h4f5 == csr_addr[11:0] ? reg_csr_1269 : _GEN_1268; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1270 = 12'h4f6 == csr_addr[11:0] ? reg_csr_1270 : _GEN_1269; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1271 = 12'h4f7 == csr_addr[11:0] ? reg_csr_1271 : _GEN_1270; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1272 = 12'h4f8 == csr_addr[11:0] ? reg_csr_1272 : _GEN_1271; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1273 = 12'h4f9 == csr_addr[11:0] ? reg_csr_1273 : _GEN_1272; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1274 = 12'h4fa == csr_addr[11:0] ? reg_csr_1274 : _GEN_1273; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1275 = 12'h4fb == csr_addr[11:0] ? reg_csr_1275 : _GEN_1274; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1276 = 12'h4fc == csr_addr[11:0] ? reg_csr_1276 : _GEN_1275; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1277 = 12'h4fd == csr_addr[11:0] ? reg_csr_1277 : _GEN_1276; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1278 = 12'h4fe == csr_addr[11:0] ? reg_csr_1278 : _GEN_1277; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1279 = 12'h4ff == csr_addr[11:0] ? reg_csr_1279 : _GEN_1278; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1280 = 12'h500 == csr_addr[11:0] ? reg_csr_1280 : _GEN_1279; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1281 = 12'h501 == csr_addr[11:0] ? reg_csr_1281 : _GEN_1280; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1282 = 12'h502 == csr_addr[11:0] ? reg_csr_1282 : _GEN_1281; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1283 = 12'h503 == csr_addr[11:0] ? reg_csr_1283 : _GEN_1282; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1284 = 12'h504 == csr_addr[11:0] ? reg_csr_1284 : _GEN_1283; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1285 = 12'h505 == csr_addr[11:0] ? reg_csr_1285 : _GEN_1284; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1286 = 12'h506 == csr_addr[11:0] ? reg_csr_1286 : _GEN_1285; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1287 = 12'h507 == csr_addr[11:0] ? reg_csr_1287 : _GEN_1286; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1288 = 12'h508 == csr_addr[11:0] ? reg_csr_1288 : _GEN_1287; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1289 = 12'h509 == csr_addr[11:0] ? reg_csr_1289 : _GEN_1288; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1290 = 12'h50a == csr_addr[11:0] ? reg_csr_1290 : _GEN_1289; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1291 = 12'h50b == csr_addr[11:0] ? reg_csr_1291 : _GEN_1290; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1292 = 12'h50c == csr_addr[11:0] ? reg_csr_1292 : _GEN_1291; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1293 = 12'h50d == csr_addr[11:0] ? reg_csr_1293 : _GEN_1292; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1294 = 12'h50e == csr_addr[11:0] ? reg_csr_1294 : _GEN_1293; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1295 = 12'h50f == csr_addr[11:0] ? reg_csr_1295 : _GEN_1294; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1296 = 12'h510 == csr_addr[11:0] ? reg_csr_1296 : _GEN_1295; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1297 = 12'h511 == csr_addr[11:0] ? reg_csr_1297 : _GEN_1296; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1298 = 12'h512 == csr_addr[11:0] ? reg_csr_1298 : _GEN_1297; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1299 = 12'h513 == csr_addr[11:0] ? reg_csr_1299 : _GEN_1298; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1300 = 12'h514 == csr_addr[11:0] ? reg_csr_1300 : _GEN_1299; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1301 = 12'h515 == csr_addr[11:0] ? reg_csr_1301 : _GEN_1300; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1302 = 12'h516 == csr_addr[11:0] ? reg_csr_1302 : _GEN_1301; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1303 = 12'h517 == csr_addr[11:0] ? reg_csr_1303 : _GEN_1302; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1304 = 12'h518 == csr_addr[11:0] ? reg_csr_1304 : _GEN_1303; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1305 = 12'h519 == csr_addr[11:0] ? reg_csr_1305 : _GEN_1304; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1306 = 12'h51a == csr_addr[11:0] ? reg_csr_1306 : _GEN_1305; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1307 = 12'h51b == csr_addr[11:0] ? reg_csr_1307 : _GEN_1306; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1308 = 12'h51c == csr_addr[11:0] ? reg_csr_1308 : _GEN_1307; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1309 = 12'h51d == csr_addr[11:0] ? reg_csr_1309 : _GEN_1308; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1310 = 12'h51e == csr_addr[11:0] ? reg_csr_1310 : _GEN_1309; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1311 = 12'h51f == csr_addr[11:0] ? reg_csr_1311 : _GEN_1310; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1312 = 12'h520 == csr_addr[11:0] ? reg_csr_1312 : _GEN_1311; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1313 = 12'h521 == csr_addr[11:0] ? reg_csr_1313 : _GEN_1312; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1314 = 12'h522 == csr_addr[11:0] ? reg_csr_1314 : _GEN_1313; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1315 = 12'h523 == csr_addr[11:0] ? reg_csr_1315 : _GEN_1314; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1316 = 12'h524 == csr_addr[11:0] ? reg_csr_1316 : _GEN_1315; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1317 = 12'h525 == csr_addr[11:0] ? reg_csr_1317 : _GEN_1316; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1318 = 12'h526 == csr_addr[11:0] ? reg_csr_1318 : _GEN_1317; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1319 = 12'h527 == csr_addr[11:0] ? reg_csr_1319 : _GEN_1318; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1320 = 12'h528 == csr_addr[11:0] ? reg_csr_1320 : _GEN_1319; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1321 = 12'h529 == csr_addr[11:0] ? reg_csr_1321 : _GEN_1320; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1322 = 12'h52a == csr_addr[11:0] ? reg_csr_1322 : _GEN_1321; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1323 = 12'h52b == csr_addr[11:0] ? reg_csr_1323 : _GEN_1322; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1324 = 12'h52c == csr_addr[11:0] ? reg_csr_1324 : _GEN_1323; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1325 = 12'h52d == csr_addr[11:0] ? reg_csr_1325 : _GEN_1324; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1326 = 12'h52e == csr_addr[11:0] ? reg_csr_1326 : _GEN_1325; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1327 = 12'h52f == csr_addr[11:0] ? reg_csr_1327 : _GEN_1326; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1328 = 12'h530 == csr_addr[11:0] ? reg_csr_1328 : _GEN_1327; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1329 = 12'h531 == csr_addr[11:0] ? reg_csr_1329 : _GEN_1328; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1330 = 12'h532 == csr_addr[11:0] ? reg_csr_1330 : _GEN_1329; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1331 = 12'h533 == csr_addr[11:0] ? reg_csr_1331 : _GEN_1330; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1332 = 12'h534 == csr_addr[11:0] ? reg_csr_1332 : _GEN_1331; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1333 = 12'h535 == csr_addr[11:0] ? reg_csr_1333 : _GEN_1332; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1334 = 12'h536 == csr_addr[11:0] ? reg_csr_1334 : _GEN_1333; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1335 = 12'h537 == csr_addr[11:0] ? reg_csr_1335 : _GEN_1334; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1336 = 12'h538 == csr_addr[11:0] ? reg_csr_1336 : _GEN_1335; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1337 = 12'h539 == csr_addr[11:0] ? reg_csr_1337 : _GEN_1336; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1338 = 12'h53a == csr_addr[11:0] ? reg_csr_1338 : _GEN_1337; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1339 = 12'h53b == csr_addr[11:0] ? reg_csr_1339 : _GEN_1338; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1340 = 12'h53c == csr_addr[11:0] ? reg_csr_1340 : _GEN_1339; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1341 = 12'h53d == csr_addr[11:0] ? reg_csr_1341 : _GEN_1340; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1342 = 12'h53e == csr_addr[11:0] ? reg_csr_1342 : _GEN_1341; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1343 = 12'h53f == csr_addr[11:0] ? reg_csr_1343 : _GEN_1342; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1344 = 12'h540 == csr_addr[11:0] ? reg_csr_1344 : _GEN_1343; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1345 = 12'h541 == csr_addr[11:0] ? reg_csr_1345 : _GEN_1344; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1346 = 12'h542 == csr_addr[11:0] ? reg_csr_1346 : _GEN_1345; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1347 = 12'h543 == csr_addr[11:0] ? reg_csr_1347 : _GEN_1346; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1348 = 12'h544 == csr_addr[11:0] ? reg_csr_1348 : _GEN_1347; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1349 = 12'h545 == csr_addr[11:0] ? reg_csr_1349 : _GEN_1348; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1350 = 12'h546 == csr_addr[11:0] ? reg_csr_1350 : _GEN_1349; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1351 = 12'h547 == csr_addr[11:0] ? reg_csr_1351 : _GEN_1350; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1352 = 12'h548 == csr_addr[11:0] ? reg_csr_1352 : _GEN_1351; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1353 = 12'h549 == csr_addr[11:0] ? reg_csr_1353 : _GEN_1352; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1354 = 12'h54a == csr_addr[11:0] ? reg_csr_1354 : _GEN_1353; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1355 = 12'h54b == csr_addr[11:0] ? reg_csr_1355 : _GEN_1354; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1356 = 12'h54c == csr_addr[11:0] ? reg_csr_1356 : _GEN_1355; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1357 = 12'h54d == csr_addr[11:0] ? reg_csr_1357 : _GEN_1356; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1358 = 12'h54e == csr_addr[11:0] ? reg_csr_1358 : _GEN_1357; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1359 = 12'h54f == csr_addr[11:0] ? reg_csr_1359 : _GEN_1358; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1360 = 12'h550 == csr_addr[11:0] ? reg_csr_1360 : _GEN_1359; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1361 = 12'h551 == csr_addr[11:0] ? reg_csr_1361 : _GEN_1360; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1362 = 12'h552 == csr_addr[11:0] ? reg_csr_1362 : _GEN_1361; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1363 = 12'h553 == csr_addr[11:0] ? reg_csr_1363 : _GEN_1362; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1364 = 12'h554 == csr_addr[11:0] ? reg_csr_1364 : _GEN_1363; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1365 = 12'h555 == csr_addr[11:0] ? reg_csr_1365 : _GEN_1364; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1366 = 12'h556 == csr_addr[11:0] ? reg_csr_1366 : _GEN_1365; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1367 = 12'h557 == csr_addr[11:0] ? reg_csr_1367 : _GEN_1366; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1368 = 12'h558 == csr_addr[11:0] ? reg_csr_1368 : _GEN_1367; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1369 = 12'h559 == csr_addr[11:0] ? reg_csr_1369 : _GEN_1368; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1370 = 12'h55a == csr_addr[11:0] ? reg_csr_1370 : _GEN_1369; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1371 = 12'h55b == csr_addr[11:0] ? reg_csr_1371 : _GEN_1370; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1372 = 12'h55c == csr_addr[11:0] ? reg_csr_1372 : _GEN_1371; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1373 = 12'h55d == csr_addr[11:0] ? reg_csr_1373 : _GEN_1372; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1374 = 12'h55e == csr_addr[11:0] ? reg_csr_1374 : _GEN_1373; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1375 = 12'h55f == csr_addr[11:0] ? reg_csr_1375 : _GEN_1374; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1376 = 12'h560 == csr_addr[11:0] ? reg_csr_1376 : _GEN_1375; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1377 = 12'h561 == csr_addr[11:0] ? reg_csr_1377 : _GEN_1376; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1378 = 12'h562 == csr_addr[11:0] ? reg_csr_1378 : _GEN_1377; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1379 = 12'h563 == csr_addr[11:0] ? reg_csr_1379 : _GEN_1378; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1380 = 12'h564 == csr_addr[11:0] ? reg_csr_1380 : _GEN_1379; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1381 = 12'h565 == csr_addr[11:0] ? reg_csr_1381 : _GEN_1380; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1382 = 12'h566 == csr_addr[11:0] ? reg_csr_1382 : _GEN_1381; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1383 = 12'h567 == csr_addr[11:0] ? reg_csr_1383 : _GEN_1382; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1384 = 12'h568 == csr_addr[11:0] ? reg_csr_1384 : _GEN_1383; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1385 = 12'h569 == csr_addr[11:0] ? reg_csr_1385 : _GEN_1384; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1386 = 12'h56a == csr_addr[11:0] ? reg_csr_1386 : _GEN_1385; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1387 = 12'h56b == csr_addr[11:0] ? reg_csr_1387 : _GEN_1386; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1388 = 12'h56c == csr_addr[11:0] ? reg_csr_1388 : _GEN_1387; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1389 = 12'h56d == csr_addr[11:0] ? reg_csr_1389 : _GEN_1388; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1390 = 12'h56e == csr_addr[11:0] ? reg_csr_1390 : _GEN_1389; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1391 = 12'h56f == csr_addr[11:0] ? reg_csr_1391 : _GEN_1390; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1392 = 12'h570 == csr_addr[11:0] ? reg_csr_1392 : _GEN_1391; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1393 = 12'h571 == csr_addr[11:0] ? reg_csr_1393 : _GEN_1392; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1394 = 12'h572 == csr_addr[11:0] ? reg_csr_1394 : _GEN_1393; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1395 = 12'h573 == csr_addr[11:0] ? reg_csr_1395 : _GEN_1394; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1396 = 12'h574 == csr_addr[11:0] ? reg_csr_1396 : _GEN_1395; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1397 = 12'h575 == csr_addr[11:0] ? reg_csr_1397 : _GEN_1396; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1398 = 12'h576 == csr_addr[11:0] ? reg_csr_1398 : _GEN_1397; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1399 = 12'h577 == csr_addr[11:0] ? reg_csr_1399 : _GEN_1398; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1400 = 12'h578 == csr_addr[11:0] ? reg_csr_1400 : _GEN_1399; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1401 = 12'h579 == csr_addr[11:0] ? reg_csr_1401 : _GEN_1400; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1402 = 12'h57a == csr_addr[11:0] ? reg_csr_1402 : _GEN_1401; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1403 = 12'h57b == csr_addr[11:0] ? reg_csr_1403 : _GEN_1402; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1404 = 12'h57c == csr_addr[11:0] ? reg_csr_1404 : _GEN_1403; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1405 = 12'h57d == csr_addr[11:0] ? reg_csr_1405 : _GEN_1404; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1406 = 12'h57e == csr_addr[11:0] ? reg_csr_1406 : _GEN_1405; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1407 = 12'h57f == csr_addr[11:0] ? reg_csr_1407 : _GEN_1406; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1408 = 12'h580 == csr_addr[11:0] ? reg_csr_1408 : _GEN_1407; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1409 = 12'h581 == csr_addr[11:0] ? reg_csr_1409 : _GEN_1408; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1410 = 12'h582 == csr_addr[11:0] ? reg_csr_1410 : _GEN_1409; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1411 = 12'h583 == csr_addr[11:0] ? reg_csr_1411 : _GEN_1410; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1412 = 12'h584 == csr_addr[11:0] ? reg_csr_1412 : _GEN_1411; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1413 = 12'h585 == csr_addr[11:0] ? reg_csr_1413 : _GEN_1412; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1414 = 12'h586 == csr_addr[11:0] ? reg_csr_1414 : _GEN_1413; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1415 = 12'h587 == csr_addr[11:0] ? reg_csr_1415 : _GEN_1414; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1416 = 12'h588 == csr_addr[11:0] ? reg_csr_1416 : _GEN_1415; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1417 = 12'h589 == csr_addr[11:0] ? reg_csr_1417 : _GEN_1416; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1418 = 12'h58a == csr_addr[11:0] ? reg_csr_1418 : _GEN_1417; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1419 = 12'h58b == csr_addr[11:0] ? reg_csr_1419 : _GEN_1418; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1420 = 12'h58c == csr_addr[11:0] ? reg_csr_1420 : _GEN_1419; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1421 = 12'h58d == csr_addr[11:0] ? reg_csr_1421 : _GEN_1420; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1422 = 12'h58e == csr_addr[11:0] ? reg_csr_1422 : _GEN_1421; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1423 = 12'h58f == csr_addr[11:0] ? reg_csr_1423 : _GEN_1422; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1424 = 12'h590 == csr_addr[11:0] ? reg_csr_1424 : _GEN_1423; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1425 = 12'h591 == csr_addr[11:0] ? reg_csr_1425 : _GEN_1424; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1426 = 12'h592 == csr_addr[11:0] ? reg_csr_1426 : _GEN_1425; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1427 = 12'h593 == csr_addr[11:0] ? reg_csr_1427 : _GEN_1426; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1428 = 12'h594 == csr_addr[11:0] ? reg_csr_1428 : _GEN_1427; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1429 = 12'h595 == csr_addr[11:0] ? reg_csr_1429 : _GEN_1428; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1430 = 12'h596 == csr_addr[11:0] ? reg_csr_1430 : _GEN_1429; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1431 = 12'h597 == csr_addr[11:0] ? reg_csr_1431 : _GEN_1430; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1432 = 12'h598 == csr_addr[11:0] ? reg_csr_1432 : _GEN_1431; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1433 = 12'h599 == csr_addr[11:0] ? reg_csr_1433 : _GEN_1432; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1434 = 12'h59a == csr_addr[11:0] ? reg_csr_1434 : _GEN_1433; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1435 = 12'h59b == csr_addr[11:0] ? reg_csr_1435 : _GEN_1434; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1436 = 12'h59c == csr_addr[11:0] ? reg_csr_1436 : _GEN_1435; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1437 = 12'h59d == csr_addr[11:0] ? reg_csr_1437 : _GEN_1436; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1438 = 12'h59e == csr_addr[11:0] ? reg_csr_1438 : _GEN_1437; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1439 = 12'h59f == csr_addr[11:0] ? reg_csr_1439 : _GEN_1438; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1440 = 12'h5a0 == csr_addr[11:0] ? reg_csr_1440 : _GEN_1439; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1441 = 12'h5a1 == csr_addr[11:0] ? reg_csr_1441 : _GEN_1440; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1442 = 12'h5a2 == csr_addr[11:0] ? reg_csr_1442 : _GEN_1441; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1443 = 12'h5a3 == csr_addr[11:0] ? reg_csr_1443 : _GEN_1442; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1444 = 12'h5a4 == csr_addr[11:0] ? reg_csr_1444 : _GEN_1443; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1445 = 12'h5a5 == csr_addr[11:0] ? reg_csr_1445 : _GEN_1444; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1446 = 12'h5a6 == csr_addr[11:0] ? reg_csr_1446 : _GEN_1445; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1447 = 12'h5a7 == csr_addr[11:0] ? reg_csr_1447 : _GEN_1446; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1448 = 12'h5a8 == csr_addr[11:0] ? reg_csr_1448 : _GEN_1447; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1449 = 12'h5a9 == csr_addr[11:0] ? reg_csr_1449 : _GEN_1448; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1450 = 12'h5aa == csr_addr[11:0] ? reg_csr_1450 : _GEN_1449; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1451 = 12'h5ab == csr_addr[11:0] ? reg_csr_1451 : _GEN_1450; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1452 = 12'h5ac == csr_addr[11:0] ? reg_csr_1452 : _GEN_1451; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1453 = 12'h5ad == csr_addr[11:0] ? reg_csr_1453 : _GEN_1452; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1454 = 12'h5ae == csr_addr[11:0] ? reg_csr_1454 : _GEN_1453; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1455 = 12'h5af == csr_addr[11:0] ? reg_csr_1455 : _GEN_1454; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1456 = 12'h5b0 == csr_addr[11:0] ? reg_csr_1456 : _GEN_1455; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1457 = 12'h5b1 == csr_addr[11:0] ? reg_csr_1457 : _GEN_1456; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1458 = 12'h5b2 == csr_addr[11:0] ? reg_csr_1458 : _GEN_1457; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1459 = 12'h5b3 == csr_addr[11:0] ? reg_csr_1459 : _GEN_1458; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1460 = 12'h5b4 == csr_addr[11:0] ? reg_csr_1460 : _GEN_1459; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1461 = 12'h5b5 == csr_addr[11:0] ? reg_csr_1461 : _GEN_1460; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1462 = 12'h5b6 == csr_addr[11:0] ? reg_csr_1462 : _GEN_1461; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1463 = 12'h5b7 == csr_addr[11:0] ? reg_csr_1463 : _GEN_1462; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1464 = 12'h5b8 == csr_addr[11:0] ? reg_csr_1464 : _GEN_1463; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1465 = 12'h5b9 == csr_addr[11:0] ? reg_csr_1465 : _GEN_1464; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1466 = 12'h5ba == csr_addr[11:0] ? reg_csr_1466 : _GEN_1465; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1467 = 12'h5bb == csr_addr[11:0] ? reg_csr_1467 : _GEN_1466; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1468 = 12'h5bc == csr_addr[11:0] ? reg_csr_1468 : _GEN_1467; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1469 = 12'h5bd == csr_addr[11:0] ? reg_csr_1469 : _GEN_1468; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1470 = 12'h5be == csr_addr[11:0] ? reg_csr_1470 : _GEN_1469; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1471 = 12'h5bf == csr_addr[11:0] ? reg_csr_1471 : _GEN_1470; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1472 = 12'h5c0 == csr_addr[11:0] ? reg_csr_1472 : _GEN_1471; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1473 = 12'h5c1 == csr_addr[11:0] ? reg_csr_1473 : _GEN_1472; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1474 = 12'h5c2 == csr_addr[11:0] ? reg_csr_1474 : _GEN_1473; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1475 = 12'h5c3 == csr_addr[11:0] ? reg_csr_1475 : _GEN_1474; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1476 = 12'h5c4 == csr_addr[11:0] ? reg_csr_1476 : _GEN_1475; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1477 = 12'h5c5 == csr_addr[11:0] ? reg_csr_1477 : _GEN_1476; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1478 = 12'h5c6 == csr_addr[11:0] ? reg_csr_1478 : _GEN_1477; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1479 = 12'h5c7 == csr_addr[11:0] ? reg_csr_1479 : _GEN_1478; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1480 = 12'h5c8 == csr_addr[11:0] ? reg_csr_1480 : _GEN_1479; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1481 = 12'h5c9 == csr_addr[11:0] ? reg_csr_1481 : _GEN_1480; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1482 = 12'h5ca == csr_addr[11:0] ? reg_csr_1482 : _GEN_1481; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1483 = 12'h5cb == csr_addr[11:0] ? reg_csr_1483 : _GEN_1482; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1484 = 12'h5cc == csr_addr[11:0] ? reg_csr_1484 : _GEN_1483; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1485 = 12'h5cd == csr_addr[11:0] ? reg_csr_1485 : _GEN_1484; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1486 = 12'h5ce == csr_addr[11:0] ? reg_csr_1486 : _GEN_1485; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1487 = 12'h5cf == csr_addr[11:0] ? reg_csr_1487 : _GEN_1486; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1488 = 12'h5d0 == csr_addr[11:0] ? reg_csr_1488 : _GEN_1487; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1489 = 12'h5d1 == csr_addr[11:0] ? reg_csr_1489 : _GEN_1488; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1490 = 12'h5d2 == csr_addr[11:0] ? reg_csr_1490 : _GEN_1489; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1491 = 12'h5d3 == csr_addr[11:0] ? reg_csr_1491 : _GEN_1490; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1492 = 12'h5d4 == csr_addr[11:0] ? reg_csr_1492 : _GEN_1491; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1493 = 12'h5d5 == csr_addr[11:0] ? reg_csr_1493 : _GEN_1492; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1494 = 12'h5d6 == csr_addr[11:0] ? reg_csr_1494 : _GEN_1493; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1495 = 12'h5d7 == csr_addr[11:0] ? reg_csr_1495 : _GEN_1494; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1496 = 12'h5d8 == csr_addr[11:0] ? reg_csr_1496 : _GEN_1495; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1497 = 12'h5d9 == csr_addr[11:0] ? reg_csr_1497 : _GEN_1496; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1498 = 12'h5da == csr_addr[11:0] ? reg_csr_1498 : _GEN_1497; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1499 = 12'h5db == csr_addr[11:0] ? reg_csr_1499 : _GEN_1498; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1500 = 12'h5dc == csr_addr[11:0] ? reg_csr_1500 : _GEN_1499; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1501 = 12'h5dd == csr_addr[11:0] ? reg_csr_1501 : _GEN_1500; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1502 = 12'h5de == csr_addr[11:0] ? reg_csr_1502 : _GEN_1501; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1503 = 12'h5df == csr_addr[11:0] ? reg_csr_1503 : _GEN_1502; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1504 = 12'h5e0 == csr_addr[11:0] ? reg_csr_1504 : _GEN_1503; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1505 = 12'h5e1 == csr_addr[11:0] ? reg_csr_1505 : _GEN_1504; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1506 = 12'h5e2 == csr_addr[11:0] ? reg_csr_1506 : _GEN_1505; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1507 = 12'h5e3 == csr_addr[11:0] ? reg_csr_1507 : _GEN_1506; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1508 = 12'h5e4 == csr_addr[11:0] ? reg_csr_1508 : _GEN_1507; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1509 = 12'h5e5 == csr_addr[11:0] ? reg_csr_1509 : _GEN_1508; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1510 = 12'h5e6 == csr_addr[11:0] ? reg_csr_1510 : _GEN_1509; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1511 = 12'h5e7 == csr_addr[11:0] ? reg_csr_1511 : _GEN_1510; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1512 = 12'h5e8 == csr_addr[11:0] ? reg_csr_1512 : _GEN_1511; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1513 = 12'h5e9 == csr_addr[11:0] ? reg_csr_1513 : _GEN_1512; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1514 = 12'h5ea == csr_addr[11:0] ? reg_csr_1514 : _GEN_1513; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1515 = 12'h5eb == csr_addr[11:0] ? reg_csr_1515 : _GEN_1514; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1516 = 12'h5ec == csr_addr[11:0] ? reg_csr_1516 : _GEN_1515; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1517 = 12'h5ed == csr_addr[11:0] ? reg_csr_1517 : _GEN_1516; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1518 = 12'h5ee == csr_addr[11:0] ? reg_csr_1518 : _GEN_1517; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1519 = 12'h5ef == csr_addr[11:0] ? reg_csr_1519 : _GEN_1518; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1520 = 12'h5f0 == csr_addr[11:0] ? reg_csr_1520 : _GEN_1519; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1521 = 12'h5f1 == csr_addr[11:0] ? reg_csr_1521 : _GEN_1520; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1522 = 12'h5f2 == csr_addr[11:0] ? reg_csr_1522 : _GEN_1521; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1523 = 12'h5f3 == csr_addr[11:0] ? reg_csr_1523 : _GEN_1522; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1524 = 12'h5f4 == csr_addr[11:0] ? reg_csr_1524 : _GEN_1523; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1525 = 12'h5f5 == csr_addr[11:0] ? reg_csr_1525 : _GEN_1524; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1526 = 12'h5f6 == csr_addr[11:0] ? reg_csr_1526 : _GEN_1525; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1527 = 12'h5f7 == csr_addr[11:0] ? reg_csr_1527 : _GEN_1526; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1528 = 12'h5f8 == csr_addr[11:0] ? reg_csr_1528 : _GEN_1527; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1529 = 12'h5f9 == csr_addr[11:0] ? reg_csr_1529 : _GEN_1528; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1530 = 12'h5fa == csr_addr[11:0] ? reg_csr_1530 : _GEN_1529; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1531 = 12'h5fb == csr_addr[11:0] ? reg_csr_1531 : _GEN_1530; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1532 = 12'h5fc == csr_addr[11:0] ? reg_csr_1532 : _GEN_1531; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1533 = 12'h5fd == csr_addr[11:0] ? reg_csr_1533 : _GEN_1532; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1534 = 12'h5fe == csr_addr[11:0] ? reg_csr_1534 : _GEN_1533; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1535 = 12'h5ff == csr_addr[11:0] ? reg_csr_1535 : _GEN_1534; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1536 = 12'h600 == csr_addr[11:0] ? reg_csr_1536 : _GEN_1535; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1537 = 12'h601 == csr_addr[11:0] ? reg_csr_1537 : _GEN_1536; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1538 = 12'h602 == csr_addr[11:0] ? reg_csr_1538 : _GEN_1537; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1539 = 12'h603 == csr_addr[11:0] ? reg_csr_1539 : _GEN_1538; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1540 = 12'h604 == csr_addr[11:0] ? reg_csr_1540 : _GEN_1539; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1541 = 12'h605 == csr_addr[11:0] ? reg_csr_1541 : _GEN_1540; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1542 = 12'h606 == csr_addr[11:0] ? reg_csr_1542 : _GEN_1541; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1543 = 12'h607 == csr_addr[11:0] ? reg_csr_1543 : _GEN_1542; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1544 = 12'h608 == csr_addr[11:0] ? reg_csr_1544 : _GEN_1543; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1545 = 12'h609 == csr_addr[11:0] ? reg_csr_1545 : _GEN_1544; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1546 = 12'h60a == csr_addr[11:0] ? reg_csr_1546 : _GEN_1545; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1547 = 12'h60b == csr_addr[11:0] ? reg_csr_1547 : _GEN_1546; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1548 = 12'h60c == csr_addr[11:0] ? reg_csr_1548 : _GEN_1547; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1549 = 12'h60d == csr_addr[11:0] ? reg_csr_1549 : _GEN_1548; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1550 = 12'h60e == csr_addr[11:0] ? reg_csr_1550 : _GEN_1549; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1551 = 12'h60f == csr_addr[11:0] ? reg_csr_1551 : _GEN_1550; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1552 = 12'h610 == csr_addr[11:0] ? reg_csr_1552 : _GEN_1551; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1553 = 12'h611 == csr_addr[11:0] ? reg_csr_1553 : _GEN_1552; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1554 = 12'h612 == csr_addr[11:0] ? reg_csr_1554 : _GEN_1553; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1555 = 12'h613 == csr_addr[11:0] ? reg_csr_1555 : _GEN_1554; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1556 = 12'h614 == csr_addr[11:0] ? reg_csr_1556 : _GEN_1555; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1557 = 12'h615 == csr_addr[11:0] ? reg_csr_1557 : _GEN_1556; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1558 = 12'h616 == csr_addr[11:0] ? reg_csr_1558 : _GEN_1557; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1559 = 12'h617 == csr_addr[11:0] ? reg_csr_1559 : _GEN_1558; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1560 = 12'h618 == csr_addr[11:0] ? reg_csr_1560 : _GEN_1559; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1561 = 12'h619 == csr_addr[11:0] ? reg_csr_1561 : _GEN_1560; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1562 = 12'h61a == csr_addr[11:0] ? reg_csr_1562 : _GEN_1561; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1563 = 12'h61b == csr_addr[11:0] ? reg_csr_1563 : _GEN_1562; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1564 = 12'h61c == csr_addr[11:0] ? reg_csr_1564 : _GEN_1563; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1565 = 12'h61d == csr_addr[11:0] ? reg_csr_1565 : _GEN_1564; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1566 = 12'h61e == csr_addr[11:0] ? reg_csr_1566 : _GEN_1565; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1567 = 12'h61f == csr_addr[11:0] ? reg_csr_1567 : _GEN_1566; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1568 = 12'h620 == csr_addr[11:0] ? reg_csr_1568 : _GEN_1567; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1569 = 12'h621 == csr_addr[11:0] ? reg_csr_1569 : _GEN_1568; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1570 = 12'h622 == csr_addr[11:0] ? reg_csr_1570 : _GEN_1569; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1571 = 12'h623 == csr_addr[11:0] ? reg_csr_1571 : _GEN_1570; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1572 = 12'h624 == csr_addr[11:0] ? reg_csr_1572 : _GEN_1571; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1573 = 12'h625 == csr_addr[11:0] ? reg_csr_1573 : _GEN_1572; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1574 = 12'h626 == csr_addr[11:0] ? reg_csr_1574 : _GEN_1573; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1575 = 12'h627 == csr_addr[11:0] ? reg_csr_1575 : _GEN_1574; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1576 = 12'h628 == csr_addr[11:0] ? reg_csr_1576 : _GEN_1575; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1577 = 12'h629 == csr_addr[11:0] ? reg_csr_1577 : _GEN_1576; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1578 = 12'h62a == csr_addr[11:0] ? reg_csr_1578 : _GEN_1577; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1579 = 12'h62b == csr_addr[11:0] ? reg_csr_1579 : _GEN_1578; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1580 = 12'h62c == csr_addr[11:0] ? reg_csr_1580 : _GEN_1579; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1581 = 12'h62d == csr_addr[11:0] ? reg_csr_1581 : _GEN_1580; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1582 = 12'h62e == csr_addr[11:0] ? reg_csr_1582 : _GEN_1581; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1583 = 12'h62f == csr_addr[11:0] ? reg_csr_1583 : _GEN_1582; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1584 = 12'h630 == csr_addr[11:0] ? reg_csr_1584 : _GEN_1583; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1585 = 12'h631 == csr_addr[11:0] ? reg_csr_1585 : _GEN_1584; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1586 = 12'h632 == csr_addr[11:0] ? reg_csr_1586 : _GEN_1585; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1587 = 12'h633 == csr_addr[11:0] ? reg_csr_1587 : _GEN_1586; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1588 = 12'h634 == csr_addr[11:0] ? reg_csr_1588 : _GEN_1587; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1589 = 12'h635 == csr_addr[11:0] ? reg_csr_1589 : _GEN_1588; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1590 = 12'h636 == csr_addr[11:0] ? reg_csr_1590 : _GEN_1589; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1591 = 12'h637 == csr_addr[11:0] ? reg_csr_1591 : _GEN_1590; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1592 = 12'h638 == csr_addr[11:0] ? reg_csr_1592 : _GEN_1591; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1593 = 12'h639 == csr_addr[11:0] ? reg_csr_1593 : _GEN_1592; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1594 = 12'h63a == csr_addr[11:0] ? reg_csr_1594 : _GEN_1593; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1595 = 12'h63b == csr_addr[11:0] ? reg_csr_1595 : _GEN_1594; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1596 = 12'h63c == csr_addr[11:0] ? reg_csr_1596 : _GEN_1595; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1597 = 12'h63d == csr_addr[11:0] ? reg_csr_1597 : _GEN_1596; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1598 = 12'h63e == csr_addr[11:0] ? reg_csr_1598 : _GEN_1597; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1599 = 12'h63f == csr_addr[11:0] ? reg_csr_1599 : _GEN_1598; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1600 = 12'h640 == csr_addr[11:0] ? reg_csr_1600 : _GEN_1599; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1601 = 12'h641 == csr_addr[11:0] ? reg_csr_1601 : _GEN_1600; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1602 = 12'h642 == csr_addr[11:0] ? reg_csr_1602 : _GEN_1601; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1603 = 12'h643 == csr_addr[11:0] ? reg_csr_1603 : _GEN_1602; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1604 = 12'h644 == csr_addr[11:0] ? reg_csr_1604 : _GEN_1603; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1605 = 12'h645 == csr_addr[11:0] ? reg_csr_1605 : _GEN_1604; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1606 = 12'h646 == csr_addr[11:0] ? reg_csr_1606 : _GEN_1605; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1607 = 12'h647 == csr_addr[11:0] ? reg_csr_1607 : _GEN_1606; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1608 = 12'h648 == csr_addr[11:0] ? reg_csr_1608 : _GEN_1607; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1609 = 12'h649 == csr_addr[11:0] ? reg_csr_1609 : _GEN_1608; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1610 = 12'h64a == csr_addr[11:0] ? reg_csr_1610 : _GEN_1609; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1611 = 12'h64b == csr_addr[11:0] ? reg_csr_1611 : _GEN_1610; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1612 = 12'h64c == csr_addr[11:0] ? reg_csr_1612 : _GEN_1611; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1613 = 12'h64d == csr_addr[11:0] ? reg_csr_1613 : _GEN_1612; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1614 = 12'h64e == csr_addr[11:0] ? reg_csr_1614 : _GEN_1613; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1615 = 12'h64f == csr_addr[11:0] ? reg_csr_1615 : _GEN_1614; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1616 = 12'h650 == csr_addr[11:0] ? reg_csr_1616 : _GEN_1615; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1617 = 12'h651 == csr_addr[11:0] ? reg_csr_1617 : _GEN_1616; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1618 = 12'h652 == csr_addr[11:0] ? reg_csr_1618 : _GEN_1617; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1619 = 12'h653 == csr_addr[11:0] ? reg_csr_1619 : _GEN_1618; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1620 = 12'h654 == csr_addr[11:0] ? reg_csr_1620 : _GEN_1619; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1621 = 12'h655 == csr_addr[11:0] ? reg_csr_1621 : _GEN_1620; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1622 = 12'h656 == csr_addr[11:0] ? reg_csr_1622 : _GEN_1621; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1623 = 12'h657 == csr_addr[11:0] ? reg_csr_1623 : _GEN_1622; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1624 = 12'h658 == csr_addr[11:0] ? reg_csr_1624 : _GEN_1623; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1625 = 12'h659 == csr_addr[11:0] ? reg_csr_1625 : _GEN_1624; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1626 = 12'h65a == csr_addr[11:0] ? reg_csr_1626 : _GEN_1625; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1627 = 12'h65b == csr_addr[11:0] ? reg_csr_1627 : _GEN_1626; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1628 = 12'h65c == csr_addr[11:0] ? reg_csr_1628 : _GEN_1627; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1629 = 12'h65d == csr_addr[11:0] ? reg_csr_1629 : _GEN_1628; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1630 = 12'h65e == csr_addr[11:0] ? reg_csr_1630 : _GEN_1629; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1631 = 12'h65f == csr_addr[11:0] ? reg_csr_1631 : _GEN_1630; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1632 = 12'h660 == csr_addr[11:0] ? reg_csr_1632 : _GEN_1631; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1633 = 12'h661 == csr_addr[11:0] ? reg_csr_1633 : _GEN_1632; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1634 = 12'h662 == csr_addr[11:0] ? reg_csr_1634 : _GEN_1633; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1635 = 12'h663 == csr_addr[11:0] ? reg_csr_1635 : _GEN_1634; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1636 = 12'h664 == csr_addr[11:0] ? reg_csr_1636 : _GEN_1635; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1637 = 12'h665 == csr_addr[11:0] ? reg_csr_1637 : _GEN_1636; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1638 = 12'h666 == csr_addr[11:0] ? reg_csr_1638 : _GEN_1637; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1639 = 12'h667 == csr_addr[11:0] ? reg_csr_1639 : _GEN_1638; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1640 = 12'h668 == csr_addr[11:0] ? reg_csr_1640 : _GEN_1639; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1641 = 12'h669 == csr_addr[11:0] ? reg_csr_1641 : _GEN_1640; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1642 = 12'h66a == csr_addr[11:0] ? reg_csr_1642 : _GEN_1641; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1643 = 12'h66b == csr_addr[11:0] ? reg_csr_1643 : _GEN_1642; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1644 = 12'h66c == csr_addr[11:0] ? reg_csr_1644 : _GEN_1643; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1645 = 12'h66d == csr_addr[11:0] ? reg_csr_1645 : _GEN_1644; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1646 = 12'h66e == csr_addr[11:0] ? reg_csr_1646 : _GEN_1645; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1647 = 12'h66f == csr_addr[11:0] ? reg_csr_1647 : _GEN_1646; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1648 = 12'h670 == csr_addr[11:0] ? reg_csr_1648 : _GEN_1647; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1649 = 12'h671 == csr_addr[11:0] ? reg_csr_1649 : _GEN_1648; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1650 = 12'h672 == csr_addr[11:0] ? reg_csr_1650 : _GEN_1649; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1651 = 12'h673 == csr_addr[11:0] ? reg_csr_1651 : _GEN_1650; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1652 = 12'h674 == csr_addr[11:0] ? reg_csr_1652 : _GEN_1651; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1653 = 12'h675 == csr_addr[11:0] ? reg_csr_1653 : _GEN_1652; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1654 = 12'h676 == csr_addr[11:0] ? reg_csr_1654 : _GEN_1653; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1655 = 12'h677 == csr_addr[11:0] ? reg_csr_1655 : _GEN_1654; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1656 = 12'h678 == csr_addr[11:0] ? reg_csr_1656 : _GEN_1655; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1657 = 12'h679 == csr_addr[11:0] ? reg_csr_1657 : _GEN_1656; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1658 = 12'h67a == csr_addr[11:0] ? reg_csr_1658 : _GEN_1657; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1659 = 12'h67b == csr_addr[11:0] ? reg_csr_1659 : _GEN_1658; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1660 = 12'h67c == csr_addr[11:0] ? reg_csr_1660 : _GEN_1659; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1661 = 12'h67d == csr_addr[11:0] ? reg_csr_1661 : _GEN_1660; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1662 = 12'h67e == csr_addr[11:0] ? reg_csr_1662 : _GEN_1661; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1663 = 12'h67f == csr_addr[11:0] ? reg_csr_1663 : _GEN_1662; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1664 = 12'h680 == csr_addr[11:0] ? reg_csr_1664 : _GEN_1663; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1665 = 12'h681 == csr_addr[11:0] ? reg_csr_1665 : _GEN_1664; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1666 = 12'h682 == csr_addr[11:0] ? reg_csr_1666 : _GEN_1665; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1667 = 12'h683 == csr_addr[11:0] ? reg_csr_1667 : _GEN_1666; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1668 = 12'h684 == csr_addr[11:0] ? reg_csr_1668 : _GEN_1667; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1669 = 12'h685 == csr_addr[11:0] ? reg_csr_1669 : _GEN_1668; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1670 = 12'h686 == csr_addr[11:0] ? reg_csr_1670 : _GEN_1669; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1671 = 12'h687 == csr_addr[11:0] ? reg_csr_1671 : _GEN_1670; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1672 = 12'h688 == csr_addr[11:0] ? reg_csr_1672 : _GEN_1671; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1673 = 12'h689 == csr_addr[11:0] ? reg_csr_1673 : _GEN_1672; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1674 = 12'h68a == csr_addr[11:0] ? reg_csr_1674 : _GEN_1673; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1675 = 12'h68b == csr_addr[11:0] ? reg_csr_1675 : _GEN_1674; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1676 = 12'h68c == csr_addr[11:0] ? reg_csr_1676 : _GEN_1675; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1677 = 12'h68d == csr_addr[11:0] ? reg_csr_1677 : _GEN_1676; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1678 = 12'h68e == csr_addr[11:0] ? reg_csr_1678 : _GEN_1677; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1679 = 12'h68f == csr_addr[11:0] ? reg_csr_1679 : _GEN_1678; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1680 = 12'h690 == csr_addr[11:0] ? reg_csr_1680 : _GEN_1679; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1681 = 12'h691 == csr_addr[11:0] ? reg_csr_1681 : _GEN_1680; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1682 = 12'h692 == csr_addr[11:0] ? reg_csr_1682 : _GEN_1681; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1683 = 12'h693 == csr_addr[11:0] ? reg_csr_1683 : _GEN_1682; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1684 = 12'h694 == csr_addr[11:0] ? reg_csr_1684 : _GEN_1683; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1685 = 12'h695 == csr_addr[11:0] ? reg_csr_1685 : _GEN_1684; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1686 = 12'h696 == csr_addr[11:0] ? reg_csr_1686 : _GEN_1685; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1687 = 12'h697 == csr_addr[11:0] ? reg_csr_1687 : _GEN_1686; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1688 = 12'h698 == csr_addr[11:0] ? reg_csr_1688 : _GEN_1687; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1689 = 12'h699 == csr_addr[11:0] ? reg_csr_1689 : _GEN_1688; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1690 = 12'h69a == csr_addr[11:0] ? reg_csr_1690 : _GEN_1689; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1691 = 12'h69b == csr_addr[11:0] ? reg_csr_1691 : _GEN_1690; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1692 = 12'h69c == csr_addr[11:0] ? reg_csr_1692 : _GEN_1691; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1693 = 12'h69d == csr_addr[11:0] ? reg_csr_1693 : _GEN_1692; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1694 = 12'h69e == csr_addr[11:0] ? reg_csr_1694 : _GEN_1693; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1695 = 12'h69f == csr_addr[11:0] ? reg_csr_1695 : _GEN_1694; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1696 = 12'h6a0 == csr_addr[11:0] ? reg_csr_1696 : _GEN_1695; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1697 = 12'h6a1 == csr_addr[11:0] ? reg_csr_1697 : _GEN_1696; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1698 = 12'h6a2 == csr_addr[11:0] ? reg_csr_1698 : _GEN_1697; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1699 = 12'h6a3 == csr_addr[11:0] ? reg_csr_1699 : _GEN_1698; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1700 = 12'h6a4 == csr_addr[11:0] ? reg_csr_1700 : _GEN_1699; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1701 = 12'h6a5 == csr_addr[11:0] ? reg_csr_1701 : _GEN_1700; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1702 = 12'h6a6 == csr_addr[11:0] ? reg_csr_1702 : _GEN_1701; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1703 = 12'h6a7 == csr_addr[11:0] ? reg_csr_1703 : _GEN_1702; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1704 = 12'h6a8 == csr_addr[11:0] ? reg_csr_1704 : _GEN_1703; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1705 = 12'h6a9 == csr_addr[11:0] ? reg_csr_1705 : _GEN_1704; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1706 = 12'h6aa == csr_addr[11:0] ? reg_csr_1706 : _GEN_1705; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1707 = 12'h6ab == csr_addr[11:0] ? reg_csr_1707 : _GEN_1706; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1708 = 12'h6ac == csr_addr[11:0] ? reg_csr_1708 : _GEN_1707; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1709 = 12'h6ad == csr_addr[11:0] ? reg_csr_1709 : _GEN_1708; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1710 = 12'h6ae == csr_addr[11:0] ? reg_csr_1710 : _GEN_1709; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1711 = 12'h6af == csr_addr[11:0] ? reg_csr_1711 : _GEN_1710; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1712 = 12'h6b0 == csr_addr[11:0] ? reg_csr_1712 : _GEN_1711; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1713 = 12'h6b1 == csr_addr[11:0] ? reg_csr_1713 : _GEN_1712; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1714 = 12'h6b2 == csr_addr[11:0] ? reg_csr_1714 : _GEN_1713; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1715 = 12'h6b3 == csr_addr[11:0] ? reg_csr_1715 : _GEN_1714; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1716 = 12'h6b4 == csr_addr[11:0] ? reg_csr_1716 : _GEN_1715; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1717 = 12'h6b5 == csr_addr[11:0] ? reg_csr_1717 : _GEN_1716; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1718 = 12'h6b6 == csr_addr[11:0] ? reg_csr_1718 : _GEN_1717; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1719 = 12'h6b7 == csr_addr[11:0] ? reg_csr_1719 : _GEN_1718; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1720 = 12'h6b8 == csr_addr[11:0] ? reg_csr_1720 : _GEN_1719; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1721 = 12'h6b9 == csr_addr[11:0] ? reg_csr_1721 : _GEN_1720; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1722 = 12'h6ba == csr_addr[11:0] ? reg_csr_1722 : _GEN_1721; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1723 = 12'h6bb == csr_addr[11:0] ? reg_csr_1723 : _GEN_1722; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1724 = 12'h6bc == csr_addr[11:0] ? reg_csr_1724 : _GEN_1723; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1725 = 12'h6bd == csr_addr[11:0] ? reg_csr_1725 : _GEN_1724; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1726 = 12'h6be == csr_addr[11:0] ? reg_csr_1726 : _GEN_1725; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1727 = 12'h6bf == csr_addr[11:0] ? reg_csr_1727 : _GEN_1726; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1728 = 12'h6c0 == csr_addr[11:0] ? reg_csr_1728 : _GEN_1727; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1729 = 12'h6c1 == csr_addr[11:0] ? reg_csr_1729 : _GEN_1728; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1730 = 12'h6c2 == csr_addr[11:0] ? reg_csr_1730 : _GEN_1729; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1731 = 12'h6c3 == csr_addr[11:0] ? reg_csr_1731 : _GEN_1730; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1732 = 12'h6c4 == csr_addr[11:0] ? reg_csr_1732 : _GEN_1731; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1733 = 12'h6c5 == csr_addr[11:0] ? reg_csr_1733 : _GEN_1732; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1734 = 12'h6c6 == csr_addr[11:0] ? reg_csr_1734 : _GEN_1733; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1735 = 12'h6c7 == csr_addr[11:0] ? reg_csr_1735 : _GEN_1734; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1736 = 12'h6c8 == csr_addr[11:0] ? reg_csr_1736 : _GEN_1735; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1737 = 12'h6c9 == csr_addr[11:0] ? reg_csr_1737 : _GEN_1736; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1738 = 12'h6ca == csr_addr[11:0] ? reg_csr_1738 : _GEN_1737; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1739 = 12'h6cb == csr_addr[11:0] ? reg_csr_1739 : _GEN_1738; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1740 = 12'h6cc == csr_addr[11:0] ? reg_csr_1740 : _GEN_1739; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1741 = 12'h6cd == csr_addr[11:0] ? reg_csr_1741 : _GEN_1740; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1742 = 12'h6ce == csr_addr[11:0] ? reg_csr_1742 : _GEN_1741; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1743 = 12'h6cf == csr_addr[11:0] ? reg_csr_1743 : _GEN_1742; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1744 = 12'h6d0 == csr_addr[11:0] ? reg_csr_1744 : _GEN_1743; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1745 = 12'h6d1 == csr_addr[11:0] ? reg_csr_1745 : _GEN_1744; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1746 = 12'h6d2 == csr_addr[11:0] ? reg_csr_1746 : _GEN_1745; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1747 = 12'h6d3 == csr_addr[11:0] ? reg_csr_1747 : _GEN_1746; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1748 = 12'h6d4 == csr_addr[11:0] ? reg_csr_1748 : _GEN_1747; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1749 = 12'h6d5 == csr_addr[11:0] ? reg_csr_1749 : _GEN_1748; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1750 = 12'h6d6 == csr_addr[11:0] ? reg_csr_1750 : _GEN_1749; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1751 = 12'h6d7 == csr_addr[11:0] ? reg_csr_1751 : _GEN_1750; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1752 = 12'h6d8 == csr_addr[11:0] ? reg_csr_1752 : _GEN_1751; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1753 = 12'h6d9 == csr_addr[11:0] ? reg_csr_1753 : _GEN_1752; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1754 = 12'h6da == csr_addr[11:0] ? reg_csr_1754 : _GEN_1753; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1755 = 12'h6db == csr_addr[11:0] ? reg_csr_1755 : _GEN_1754; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1756 = 12'h6dc == csr_addr[11:0] ? reg_csr_1756 : _GEN_1755; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1757 = 12'h6dd == csr_addr[11:0] ? reg_csr_1757 : _GEN_1756; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1758 = 12'h6de == csr_addr[11:0] ? reg_csr_1758 : _GEN_1757; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1759 = 12'h6df == csr_addr[11:0] ? reg_csr_1759 : _GEN_1758; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1760 = 12'h6e0 == csr_addr[11:0] ? reg_csr_1760 : _GEN_1759; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1761 = 12'h6e1 == csr_addr[11:0] ? reg_csr_1761 : _GEN_1760; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1762 = 12'h6e2 == csr_addr[11:0] ? reg_csr_1762 : _GEN_1761; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1763 = 12'h6e3 == csr_addr[11:0] ? reg_csr_1763 : _GEN_1762; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1764 = 12'h6e4 == csr_addr[11:0] ? reg_csr_1764 : _GEN_1763; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1765 = 12'h6e5 == csr_addr[11:0] ? reg_csr_1765 : _GEN_1764; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1766 = 12'h6e6 == csr_addr[11:0] ? reg_csr_1766 : _GEN_1765; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1767 = 12'h6e7 == csr_addr[11:0] ? reg_csr_1767 : _GEN_1766; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1768 = 12'h6e8 == csr_addr[11:0] ? reg_csr_1768 : _GEN_1767; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1769 = 12'h6e9 == csr_addr[11:0] ? reg_csr_1769 : _GEN_1768; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1770 = 12'h6ea == csr_addr[11:0] ? reg_csr_1770 : _GEN_1769; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1771 = 12'h6eb == csr_addr[11:0] ? reg_csr_1771 : _GEN_1770; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1772 = 12'h6ec == csr_addr[11:0] ? reg_csr_1772 : _GEN_1771; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1773 = 12'h6ed == csr_addr[11:0] ? reg_csr_1773 : _GEN_1772; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1774 = 12'h6ee == csr_addr[11:0] ? reg_csr_1774 : _GEN_1773; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1775 = 12'h6ef == csr_addr[11:0] ? reg_csr_1775 : _GEN_1774; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1776 = 12'h6f0 == csr_addr[11:0] ? reg_csr_1776 : _GEN_1775; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1777 = 12'h6f1 == csr_addr[11:0] ? reg_csr_1777 : _GEN_1776; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1778 = 12'h6f2 == csr_addr[11:0] ? reg_csr_1778 : _GEN_1777; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1779 = 12'h6f3 == csr_addr[11:0] ? reg_csr_1779 : _GEN_1778; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1780 = 12'h6f4 == csr_addr[11:0] ? reg_csr_1780 : _GEN_1779; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1781 = 12'h6f5 == csr_addr[11:0] ? reg_csr_1781 : _GEN_1780; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1782 = 12'h6f6 == csr_addr[11:0] ? reg_csr_1782 : _GEN_1781; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1783 = 12'h6f7 == csr_addr[11:0] ? reg_csr_1783 : _GEN_1782; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1784 = 12'h6f8 == csr_addr[11:0] ? reg_csr_1784 : _GEN_1783; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1785 = 12'h6f9 == csr_addr[11:0] ? reg_csr_1785 : _GEN_1784; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1786 = 12'h6fa == csr_addr[11:0] ? reg_csr_1786 : _GEN_1785; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1787 = 12'h6fb == csr_addr[11:0] ? reg_csr_1787 : _GEN_1786; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1788 = 12'h6fc == csr_addr[11:0] ? reg_csr_1788 : _GEN_1787; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1789 = 12'h6fd == csr_addr[11:0] ? reg_csr_1789 : _GEN_1788; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1790 = 12'h6fe == csr_addr[11:0] ? reg_csr_1790 : _GEN_1789; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1791 = 12'h6ff == csr_addr[11:0] ? reg_csr_1791 : _GEN_1790; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1792 = 12'h700 == csr_addr[11:0] ? reg_csr_1792 : _GEN_1791; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1793 = 12'h701 == csr_addr[11:0] ? reg_csr_1793 : _GEN_1792; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1794 = 12'h702 == csr_addr[11:0] ? reg_csr_1794 : _GEN_1793; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1795 = 12'h703 == csr_addr[11:0] ? reg_csr_1795 : _GEN_1794; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1796 = 12'h704 == csr_addr[11:0] ? reg_csr_1796 : _GEN_1795; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1797 = 12'h705 == csr_addr[11:0] ? reg_csr_1797 : _GEN_1796; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1798 = 12'h706 == csr_addr[11:0] ? reg_csr_1798 : _GEN_1797; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1799 = 12'h707 == csr_addr[11:0] ? reg_csr_1799 : _GEN_1798; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1800 = 12'h708 == csr_addr[11:0] ? reg_csr_1800 : _GEN_1799; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1801 = 12'h709 == csr_addr[11:0] ? reg_csr_1801 : _GEN_1800; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1802 = 12'h70a == csr_addr[11:0] ? reg_csr_1802 : _GEN_1801; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1803 = 12'h70b == csr_addr[11:0] ? reg_csr_1803 : _GEN_1802; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1804 = 12'h70c == csr_addr[11:0] ? reg_csr_1804 : _GEN_1803; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1805 = 12'h70d == csr_addr[11:0] ? reg_csr_1805 : _GEN_1804; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1806 = 12'h70e == csr_addr[11:0] ? reg_csr_1806 : _GEN_1805; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1807 = 12'h70f == csr_addr[11:0] ? reg_csr_1807 : _GEN_1806; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1808 = 12'h710 == csr_addr[11:0] ? reg_csr_1808 : _GEN_1807; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1809 = 12'h711 == csr_addr[11:0] ? reg_csr_1809 : _GEN_1808; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1810 = 12'h712 == csr_addr[11:0] ? reg_csr_1810 : _GEN_1809; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1811 = 12'h713 == csr_addr[11:0] ? reg_csr_1811 : _GEN_1810; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1812 = 12'h714 == csr_addr[11:0] ? reg_csr_1812 : _GEN_1811; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1813 = 12'h715 == csr_addr[11:0] ? reg_csr_1813 : _GEN_1812; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1814 = 12'h716 == csr_addr[11:0] ? reg_csr_1814 : _GEN_1813; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1815 = 12'h717 == csr_addr[11:0] ? reg_csr_1815 : _GEN_1814; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1816 = 12'h718 == csr_addr[11:0] ? reg_csr_1816 : _GEN_1815; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1817 = 12'h719 == csr_addr[11:0] ? reg_csr_1817 : _GEN_1816; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1818 = 12'h71a == csr_addr[11:0] ? reg_csr_1818 : _GEN_1817; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1819 = 12'h71b == csr_addr[11:0] ? reg_csr_1819 : _GEN_1818; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1820 = 12'h71c == csr_addr[11:0] ? reg_csr_1820 : _GEN_1819; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1821 = 12'h71d == csr_addr[11:0] ? reg_csr_1821 : _GEN_1820; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1822 = 12'h71e == csr_addr[11:0] ? reg_csr_1822 : _GEN_1821; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1823 = 12'h71f == csr_addr[11:0] ? reg_csr_1823 : _GEN_1822; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1824 = 12'h720 == csr_addr[11:0] ? reg_csr_1824 : _GEN_1823; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1825 = 12'h721 == csr_addr[11:0] ? reg_csr_1825 : _GEN_1824; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1826 = 12'h722 == csr_addr[11:0] ? reg_csr_1826 : _GEN_1825; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1827 = 12'h723 == csr_addr[11:0] ? reg_csr_1827 : _GEN_1826; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1828 = 12'h724 == csr_addr[11:0] ? reg_csr_1828 : _GEN_1827; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1829 = 12'h725 == csr_addr[11:0] ? reg_csr_1829 : _GEN_1828; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1830 = 12'h726 == csr_addr[11:0] ? reg_csr_1830 : _GEN_1829; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1831 = 12'h727 == csr_addr[11:0] ? reg_csr_1831 : _GEN_1830; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1832 = 12'h728 == csr_addr[11:0] ? reg_csr_1832 : _GEN_1831; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1833 = 12'h729 == csr_addr[11:0] ? reg_csr_1833 : _GEN_1832; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1834 = 12'h72a == csr_addr[11:0] ? reg_csr_1834 : _GEN_1833; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1835 = 12'h72b == csr_addr[11:0] ? reg_csr_1835 : _GEN_1834; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1836 = 12'h72c == csr_addr[11:0] ? reg_csr_1836 : _GEN_1835; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1837 = 12'h72d == csr_addr[11:0] ? reg_csr_1837 : _GEN_1836; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1838 = 12'h72e == csr_addr[11:0] ? reg_csr_1838 : _GEN_1837; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1839 = 12'h72f == csr_addr[11:0] ? reg_csr_1839 : _GEN_1838; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1840 = 12'h730 == csr_addr[11:0] ? reg_csr_1840 : _GEN_1839; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1841 = 12'h731 == csr_addr[11:0] ? reg_csr_1841 : _GEN_1840; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1842 = 12'h732 == csr_addr[11:0] ? reg_csr_1842 : _GEN_1841; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1843 = 12'h733 == csr_addr[11:0] ? reg_csr_1843 : _GEN_1842; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1844 = 12'h734 == csr_addr[11:0] ? reg_csr_1844 : _GEN_1843; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1845 = 12'h735 == csr_addr[11:0] ? reg_csr_1845 : _GEN_1844; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1846 = 12'h736 == csr_addr[11:0] ? reg_csr_1846 : _GEN_1845; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1847 = 12'h737 == csr_addr[11:0] ? reg_csr_1847 : _GEN_1846; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1848 = 12'h738 == csr_addr[11:0] ? reg_csr_1848 : _GEN_1847; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1849 = 12'h739 == csr_addr[11:0] ? reg_csr_1849 : _GEN_1848; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1850 = 12'h73a == csr_addr[11:0] ? reg_csr_1850 : _GEN_1849; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1851 = 12'h73b == csr_addr[11:0] ? reg_csr_1851 : _GEN_1850; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1852 = 12'h73c == csr_addr[11:0] ? reg_csr_1852 : _GEN_1851; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1853 = 12'h73d == csr_addr[11:0] ? reg_csr_1853 : _GEN_1852; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1854 = 12'h73e == csr_addr[11:0] ? reg_csr_1854 : _GEN_1853; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1855 = 12'h73f == csr_addr[11:0] ? reg_csr_1855 : _GEN_1854; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1856 = 12'h740 == csr_addr[11:0] ? reg_csr_1856 : _GEN_1855; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1857 = 12'h741 == csr_addr[11:0] ? reg_csr_1857 : _GEN_1856; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1858 = 12'h742 == csr_addr[11:0] ? reg_csr_1858 : _GEN_1857; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1859 = 12'h743 == csr_addr[11:0] ? reg_csr_1859 : _GEN_1858; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1860 = 12'h744 == csr_addr[11:0] ? reg_csr_1860 : _GEN_1859; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1861 = 12'h745 == csr_addr[11:0] ? reg_csr_1861 : _GEN_1860; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1862 = 12'h746 == csr_addr[11:0] ? reg_csr_1862 : _GEN_1861; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1863 = 12'h747 == csr_addr[11:0] ? reg_csr_1863 : _GEN_1862; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1864 = 12'h748 == csr_addr[11:0] ? reg_csr_1864 : _GEN_1863; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1865 = 12'h749 == csr_addr[11:0] ? reg_csr_1865 : _GEN_1864; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1866 = 12'h74a == csr_addr[11:0] ? reg_csr_1866 : _GEN_1865; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1867 = 12'h74b == csr_addr[11:0] ? reg_csr_1867 : _GEN_1866; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1868 = 12'h74c == csr_addr[11:0] ? reg_csr_1868 : _GEN_1867; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1869 = 12'h74d == csr_addr[11:0] ? reg_csr_1869 : _GEN_1868; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1870 = 12'h74e == csr_addr[11:0] ? reg_csr_1870 : _GEN_1869; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1871 = 12'h74f == csr_addr[11:0] ? reg_csr_1871 : _GEN_1870; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1872 = 12'h750 == csr_addr[11:0] ? reg_csr_1872 : _GEN_1871; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1873 = 12'h751 == csr_addr[11:0] ? reg_csr_1873 : _GEN_1872; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1874 = 12'h752 == csr_addr[11:0] ? reg_csr_1874 : _GEN_1873; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1875 = 12'h753 == csr_addr[11:0] ? reg_csr_1875 : _GEN_1874; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1876 = 12'h754 == csr_addr[11:0] ? reg_csr_1876 : _GEN_1875; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1877 = 12'h755 == csr_addr[11:0] ? reg_csr_1877 : _GEN_1876; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1878 = 12'h756 == csr_addr[11:0] ? reg_csr_1878 : _GEN_1877; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1879 = 12'h757 == csr_addr[11:0] ? reg_csr_1879 : _GEN_1878; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1880 = 12'h758 == csr_addr[11:0] ? reg_csr_1880 : _GEN_1879; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1881 = 12'h759 == csr_addr[11:0] ? reg_csr_1881 : _GEN_1880; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1882 = 12'h75a == csr_addr[11:0] ? reg_csr_1882 : _GEN_1881; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1883 = 12'h75b == csr_addr[11:0] ? reg_csr_1883 : _GEN_1882; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1884 = 12'h75c == csr_addr[11:0] ? reg_csr_1884 : _GEN_1883; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1885 = 12'h75d == csr_addr[11:0] ? reg_csr_1885 : _GEN_1884; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1886 = 12'h75e == csr_addr[11:0] ? reg_csr_1886 : _GEN_1885; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1887 = 12'h75f == csr_addr[11:0] ? reg_csr_1887 : _GEN_1886; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1888 = 12'h760 == csr_addr[11:0] ? reg_csr_1888 : _GEN_1887; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1889 = 12'h761 == csr_addr[11:0] ? reg_csr_1889 : _GEN_1888; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1890 = 12'h762 == csr_addr[11:0] ? reg_csr_1890 : _GEN_1889; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1891 = 12'h763 == csr_addr[11:0] ? reg_csr_1891 : _GEN_1890; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1892 = 12'h764 == csr_addr[11:0] ? reg_csr_1892 : _GEN_1891; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1893 = 12'h765 == csr_addr[11:0] ? reg_csr_1893 : _GEN_1892; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1894 = 12'h766 == csr_addr[11:0] ? reg_csr_1894 : _GEN_1893; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1895 = 12'h767 == csr_addr[11:0] ? reg_csr_1895 : _GEN_1894; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1896 = 12'h768 == csr_addr[11:0] ? reg_csr_1896 : _GEN_1895; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1897 = 12'h769 == csr_addr[11:0] ? reg_csr_1897 : _GEN_1896; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1898 = 12'h76a == csr_addr[11:0] ? reg_csr_1898 : _GEN_1897; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1899 = 12'h76b == csr_addr[11:0] ? reg_csr_1899 : _GEN_1898; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1900 = 12'h76c == csr_addr[11:0] ? reg_csr_1900 : _GEN_1899; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1901 = 12'h76d == csr_addr[11:0] ? reg_csr_1901 : _GEN_1900; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1902 = 12'h76e == csr_addr[11:0] ? reg_csr_1902 : _GEN_1901; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1903 = 12'h76f == csr_addr[11:0] ? reg_csr_1903 : _GEN_1902; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1904 = 12'h770 == csr_addr[11:0] ? reg_csr_1904 : _GEN_1903; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1905 = 12'h771 == csr_addr[11:0] ? reg_csr_1905 : _GEN_1904; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1906 = 12'h772 == csr_addr[11:0] ? reg_csr_1906 : _GEN_1905; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1907 = 12'h773 == csr_addr[11:0] ? reg_csr_1907 : _GEN_1906; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1908 = 12'h774 == csr_addr[11:0] ? reg_csr_1908 : _GEN_1907; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1909 = 12'h775 == csr_addr[11:0] ? reg_csr_1909 : _GEN_1908; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1910 = 12'h776 == csr_addr[11:0] ? reg_csr_1910 : _GEN_1909; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1911 = 12'h777 == csr_addr[11:0] ? reg_csr_1911 : _GEN_1910; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1912 = 12'h778 == csr_addr[11:0] ? reg_csr_1912 : _GEN_1911; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1913 = 12'h779 == csr_addr[11:0] ? reg_csr_1913 : _GEN_1912; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1914 = 12'h77a == csr_addr[11:0] ? reg_csr_1914 : _GEN_1913; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1915 = 12'h77b == csr_addr[11:0] ? reg_csr_1915 : _GEN_1914; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1916 = 12'h77c == csr_addr[11:0] ? reg_csr_1916 : _GEN_1915; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1917 = 12'h77d == csr_addr[11:0] ? reg_csr_1917 : _GEN_1916; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1918 = 12'h77e == csr_addr[11:0] ? reg_csr_1918 : _GEN_1917; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1919 = 12'h77f == csr_addr[11:0] ? reg_csr_1919 : _GEN_1918; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1920 = 12'h780 == csr_addr[11:0] ? reg_csr_1920 : _GEN_1919; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1921 = 12'h781 == csr_addr[11:0] ? reg_csr_1921 : _GEN_1920; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1922 = 12'h782 == csr_addr[11:0] ? reg_csr_1922 : _GEN_1921; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1923 = 12'h783 == csr_addr[11:0] ? reg_csr_1923 : _GEN_1922; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1924 = 12'h784 == csr_addr[11:0] ? reg_csr_1924 : _GEN_1923; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1925 = 12'h785 == csr_addr[11:0] ? reg_csr_1925 : _GEN_1924; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1926 = 12'h786 == csr_addr[11:0] ? reg_csr_1926 : _GEN_1925; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1927 = 12'h787 == csr_addr[11:0] ? reg_csr_1927 : _GEN_1926; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1928 = 12'h788 == csr_addr[11:0] ? reg_csr_1928 : _GEN_1927; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1929 = 12'h789 == csr_addr[11:0] ? reg_csr_1929 : _GEN_1928; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1930 = 12'h78a == csr_addr[11:0] ? reg_csr_1930 : _GEN_1929; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1931 = 12'h78b == csr_addr[11:0] ? reg_csr_1931 : _GEN_1930; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1932 = 12'h78c == csr_addr[11:0] ? reg_csr_1932 : _GEN_1931; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1933 = 12'h78d == csr_addr[11:0] ? reg_csr_1933 : _GEN_1932; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1934 = 12'h78e == csr_addr[11:0] ? reg_csr_1934 : _GEN_1933; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1935 = 12'h78f == csr_addr[11:0] ? reg_csr_1935 : _GEN_1934; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1936 = 12'h790 == csr_addr[11:0] ? reg_csr_1936 : _GEN_1935; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1937 = 12'h791 == csr_addr[11:0] ? reg_csr_1937 : _GEN_1936; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1938 = 12'h792 == csr_addr[11:0] ? reg_csr_1938 : _GEN_1937; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1939 = 12'h793 == csr_addr[11:0] ? reg_csr_1939 : _GEN_1938; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1940 = 12'h794 == csr_addr[11:0] ? reg_csr_1940 : _GEN_1939; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1941 = 12'h795 == csr_addr[11:0] ? reg_csr_1941 : _GEN_1940; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1942 = 12'h796 == csr_addr[11:0] ? reg_csr_1942 : _GEN_1941; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1943 = 12'h797 == csr_addr[11:0] ? reg_csr_1943 : _GEN_1942; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1944 = 12'h798 == csr_addr[11:0] ? reg_csr_1944 : _GEN_1943; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1945 = 12'h799 == csr_addr[11:0] ? reg_csr_1945 : _GEN_1944; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1946 = 12'h79a == csr_addr[11:0] ? reg_csr_1946 : _GEN_1945; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1947 = 12'h79b == csr_addr[11:0] ? reg_csr_1947 : _GEN_1946; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1948 = 12'h79c == csr_addr[11:0] ? reg_csr_1948 : _GEN_1947; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1949 = 12'h79d == csr_addr[11:0] ? reg_csr_1949 : _GEN_1948; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1950 = 12'h79e == csr_addr[11:0] ? reg_csr_1950 : _GEN_1949; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1951 = 12'h79f == csr_addr[11:0] ? reg_csr_1951 : _GEN_1950; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1952 = 12'h7a0 == csr_addr[11:0] ? reg_csr_1952 : _GEN_1951; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1953 = 12'h7a1 == csr_addr[11:0] ? reg_csr_1953 : _GEN_1952; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1954 = 12'h7a2 == csr_addr[11:0] ? reg_csr_1954 : _GEN_1953; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1955 = 12'h7a3 == csr_addr[11:0] ? reg_csr_1955 : _GEN_1954; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1956 = 12'h7a4 == csr_addr[11:0] ? reg_csr_1956 : _GEN_1955; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1957 = 12'h7a5 == csr_addr[11:0] ? reg_csr_1957 : _GEN_1956; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1958 = 12'h7a6 == csr_addr[11:0] ? reg_csr_1958 : _GEN_1957; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1959 = 12'h7a7 == csr_addr[11:0] ? reg_csr_1959 : _GEN_1958; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1960 = 12'h7a8 == csr_addr[11:0] ? reg_csr_1960 : _GEN_1959; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1961 = 12'h7a9 == csr_addr[11:0] ? reg_csr_1961 : _GEN_1960; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1962 = 12'h7aa == csr_addr[11:0] ? reg_csr_1962 : _GEN_1961; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1963 = 12'h7ab == csr_addr[11:0] ? reg_csr_1963 : _GEN_1962; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1964 = 12'h7ac == csr_addr[11:0] ? reg_csr_1964 : _GEN_1963; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1965 = 12'h7ad == csr_addr[11:0] ? reg_csr_1965 : _GEN_1964; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1966 = 12'h7ae == csr_addr[11:0] ? reg_csr_1966 : _GEN_1965; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1967 = 12'h7af == csr_addr[11:0] ? reg_csr_1967 : _GEN_1966; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1968 = 12'h7b0 == csr_addr[11:0] ? reg_csr_1968 : _GEN_1967; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1969 = 12'h7b1 == csr_addr[11:0] ? reg_csr_1969 : _GEN_1968; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1970 = 12'h7b2 == csr_addr[11:0] ? reg_csr_1970 : _GEN_1969; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1971 = 12'h7b3 == csr_addr[11:0] ? reg_csr_1971 : _GEN_1970; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1972 = 12'h7b4 == csr_addr[11:0] ? reg_csr_1972 : _GEN_1971; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1973 = 12'h7b5 == csr_addr[11:0] ? reg_csr_1973 : _GEN_1972; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1974 = 12'h7b6 == csr_addr[11:0] ? reg_csr_1974 : _GEN_1973; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1975 = 12'h7b7 == csr_addr[11:0] ? reg_csr_1975 : _GEN_1974; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1976 = 12'h7b8 == csr_addr[11:0] ? reg_csr_1976 : _GEN_1975; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1977 = 12'h7b9 == csr_addr[11:0] ? reg_csr_1977 : _GEN_1976; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1978 = 12'h7ba == csr_addr[11:0] ? reg_csr_1978 : _GEN_1977; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1979 = 12'h7bb == csr_addr[11:0] ? reg_csr_1979 : _GEN_1978; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1980 = 12'h7bc == csr_addr[11:0] ? reg_csr_1980 : _GEN_1979; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1981 = 12'h7bd == csr_addr[11:0] ? reg_csr_1981 : _GEN_1980; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1982 = 12'h7be == csr_addr[11:0] ? reg_csr_1982 : _GEN_1981; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1983 = 12'h7bf == csr_addr[11:0] ? reg_csr_1983 : _GEN_1982; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1984 = 12'h7c0 == csr_addr[11:0] ? reg_csr_1984 : _GEN_1983; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1985 = 12'h7c1 == csr_addr[11:0] ? reg_csr_1985 : _GEN_1984; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1986 = 12'h7c2 == csr_addr[11:0] ? reg_csr_1986 : _GEN_1985; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1987 = 12'h7c3 == csr_addr[11:0] ? reg_csr_1987 : _GEN_1986; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1988 = 12'h7c4 == csr_addr[11:0] ? reg_csr_1988 : _GEN_1987; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1989 = 12'h7c5 == csr_addr[11:0] ? reg_csr_1989 : _GEN_1988; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1990 = 12'h7c6 == csr_addr[11:0] ? reg_csr_1990 : _GEN_1989; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1991 = 12'h7c7 == csr_addr[11:0] ? reg_csr_1991 : _GEN_1990; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1992 = 12'h7c8 == csr_addr[11:0] ? reg_csr_1992 : _GEN_1991; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1993 = 12'h7c9 == csr_addr[11:0] ? reg_csr_1993 : _GEN_1992; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1994 = 12'h7ca == csr_addr[11:0] ? reg_csr_1994 : _GEN_1993; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1995 = 12'h7cb == csr_addr[11:0] ? reg_csr_1995 : _GEN_1994; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1996 = 12'h7cc == csr_addr[11:0] ? reg_csr_1996 : _GEN_1995; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1997 = 12'h7cd == csr_addr[11:0] ? reg_csr_1997 : _GEN_1996; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1998 = 12'h7ce == csr_addr[11:0] ? reg_csr_1998 : _GEN_1997; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_1999 = 12'h7cf == csr_addr[11:0] ? reg_csr_1999 : _GEN_1998; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2000 = 12'h7d0 == csr_addr[11:0] ? reg_csr_2000 : _GEN_1999; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2001 = 12'h7d1 == csr_addr[11:0] ? reg_csr_2001 : _GEN_2000; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2002 = 12'h7d2 == csr_addr[11:0] ? reg_csr_2002 : _GEN_2001; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2003 = 12'h7d3 == csr_addr[11:0] ? reg_csr_2003 : _GEN_2002; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2004 = 12'h7d4 == csr_addr[11:0] ? reg_csr_2004 : _GEN_2003; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2005 = 12'h7d5 == csr_addr[11:0] ? reg_csr_2005 : _GEN_2004; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2006 = 12'h7d6 == csr_addr[11:0] ? reg_csr_2006 : _GEN_2005; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2007 = 12'h7d7 == csr_addr[11:0] ? reg_csr_2007 : _GEN_2006; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2008 = 12'h7d8 == csr_addr[11:0] ? reg_csr_2008 : _GEN_2007; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2009 = 12'h7d9 == csr_addr[11:0] ? reg_csr_2009 : _GEN_2008; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2010 = 12'h7da == csr_addr[11:0] ? reg_csr_2010 : _GEN_2009; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2011 = 12'h7db == csr_addr[11:0] ? reg_csr_2011 : _GEN_2010; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2012 = 12'h7dc == csr_addr[11:0] ? reg_csr_2012 : _GEN_2011; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2013 = 12'h7dd == csr_addr[11:0] ? reg_csr_2013 : _GEN_2012; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2014 = 12'h7de == csr_addr[11:0] ? reg_csr_2014 : _GEN_2013; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2015 = 12'h7df == csr_addr[11:0] ? reg_csr_2015 : _GEN_2014; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2016 = 12'h7e0 == csr_addr[11:0] ? reg_csr_2016 : _GEN_2015; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2017 = 12'h7e1 == csr_addr[11:0] ? reg_csr_2017 : _GEN_2016; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2018 = 12'h7e2 == csr_addr[11:0] ? reg_csr_2018 : _GEN_2017; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2019 = 12'h7e3 == csr_addr[11:0] ? reg_csr_2019 : _GEN_2018; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2020 = 12'h7e4 == csr_addr[11:0] ? reg_csr_2020 : _GEN_2019; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2021 = 12'h7e5 == csr_addr[11:0] ? reg_csr_2021 : _GEN_2020; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2022 = 12'h7e6 == csr_addr[11:0] ? reg_csr_2022 : _GEN_2021; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2023 = 12'h7e7 == csr_addr[11:0] ? reg_csr_2023 : _GEN_2022; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2024 = 12'h7e8 == csr_addr[11:0] ? reg_csr_2024 : _GEN_2023; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2025 = 12'h7e9 == csr_addr[11:0] ? reg_csr_2025 : _GEN_2024; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2026 = 12'h7ea == csr_addr[11:0] ? reg_csr_2026 : _GEN_2025; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2027 = 12'h7eb == csr_addr[11:0] ? reg_csr_2027 : _GEN_2026; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2028 = 12'h7ec == csr_addr[11:0] ? reg_csr_2028 : _GEN_2027; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2029 = 12'h7ed == csr_addr[11:0] ? reg_csr_2029 : _GEN_2028; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2030 = 12'h7ee == csr_addr[11:0] ? reg_csr_2030 : _GEN_2029; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2031 = 12'h7ef == csr_addr[11:0] ? reg_csr_2031 : _GEN_2030; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2032 = 12'h7f0 == csr_addr[11:0] ? reg_csr_2032 : _GEN_2031; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2033 = 12'h7f1 == csr_addr[11:0] ? reg_csr_2033 : _GEN_2032; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2034 = 12'h7f2 == csr_addr[11:0] ? reg_csr_2034 : _GEN_2033; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2035 = 12'h7f3 == csr_addr[11:0] ? reg_csr_2035 : _GEN_2034; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2036 = 12'h7f4 == csr_addr[11:0] ? reg_csr_2036 : _GEN_2035; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2037 = 12'h7f5 == csr_addr[11:0] ? reg_csr_2037 : _GEN_2036; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2038 = 12'h7f6 == csr_addr[11:0] ? reg_csr_2038 : _GEN_2037; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2039 = 12'h7f7 == csr_addr[11:0] ? reg_csr_2039 : _GEN_2038; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2040 = 12'h7f8 == csr_addr[11:0] ? reg_csr_2040 : _GEN_2039; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2041 = 12'h7f9 == csr_addr[11:0] ? reg_csr_2041 : _GEN_2040; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2042 = 12'h7fa == csr_addr[11:0] ? reg_csr_2042 : _GEN_2041; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2043 = 12'h7fb == csr_addr[11:0] ? reg_csr_2043 : _GEN_2042; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2044 = 12'h7fc == csr_addr[11:0] ? reg_csr_2044 : _GEN_2043; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2045 = 12'h7fd == csr_addr[11:0] ? reg_csr_2045 : _GEN_2044; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2046 = 12'h7fe == csr_addr[11:0] ? reg_csr_2046 : _GEN_2045; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2047 = 12'h7ff == csr_addr[11:0] ? reg_csr_2047 : _GEN_2046; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2048 = 12'h800 == csr_addr[11:0] ? reg_csr_2048 : _GEN_2047; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2049 = 12'h801 == csr_addr[11:0] ? reg_csr_2049 : _GEN_2048; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2050 = 12'h802 == csr_addr[11:0] ? reg_csr_2050 : _GEN_2049; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2051 = 12'h803 == csr_addr[11:0] ? reg_csr_2051 : _GEN_2050; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2052 = 12'h804 == csr_addr[11:0] ? reg_csr_2052 : _GEN_2051; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2053 = 12'h805 == csr_addr[11:0] ? reg_csr_2053 : _GEN_2052; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2054 = 12'h806 == csr_addr[11:0] ? reg_csr_2054 : _GEN_2053; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2055 = 12'h807 == csr_addr[11:0] ? reg_csr_2055 : _GEN_2054; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2056 = 12'h808 == csr_addr[11:0] ? reg_csr_2056 : _GEN_2055; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2057 = 12'h809 == csr_addr[11:0] ? reg_csr_2057 : _GEN_2056; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2058 = 12'h80a == csr_addr[11:0] ? reg_csr_2058 : _GEN_2057; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2059 = 12'h80b == csr_addr[11:0] ? reg_csr_2059 : _GEN_2058; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2060 = 12'h80c == csr_addr[11:0] ? reg_csr_2060 : _GEN_2059; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2061 = 12'h80d == csr_addr[11:0] ? reg_csr_2061 : _GEN_2060; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2062 = 12'h80e == csr_addr[11:0] ? reg_csr_2062 : _GEN_2061; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2063 = 12'h80f == csr_addr[11:0] ? reg_csr_2063 : _GEN_2062; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2064 = 12'h810 == csr_addr[11:0] ? reg_csr_2064 : _GEN_2063; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2065 = 12'h811 == csr_addr[11:0] ? reg_csr_2065 : _GEN_2064; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2066 = 12'h812 == csr_addr[11:0] ? reg_csr_2066 : _GEN_2065; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2067 = 12'h813 == csr_addr[11:0] ? reg_csr_2067 : _GEN_2066; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2068 = 12'h814 == csr_addr[11:0] ? reg_csr_2068 : _GEN_2067; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2069 = 12'h815 == csr_addr[11:0] ? reg_csr_2069 : _GEN_2068; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2070 = 12'h816 == csr_addr[11:0] ? reg_csr_2070 : _GEN_2069; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2071 = 12'h817 == csr_addr[11:0] ? reg_csr_2071 : _GEN_2070; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2072 = 12'h818 == csr_addr[11:0] ? reg_csr_2072 : _GEN_2071; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2073 = 12'h819 == csr_addr[11:0] ? reg_csr_2073 : _GEN_2072; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2074 = 12'h81a == csr_addr[11:0] ? reg_csr_2074 : _GEN_2073; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2075 = 12'h81b == csr_addr[11:0] ? reg_csr_2075 : _GEN_2074; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2076 = 12'h81c == csr_addr[11:0] ? reg_csr_2076 : _GEN_2075; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2077 = 12'h81d == csr_addr[11:0] ? reg_csr_2077 : _GEN_2076; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2078 = 12'h81e == csr_addr[11:0] ? reg_csr_2078 : _GEN_2077; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2079 = 12'h81f == csr_addr[11:0] ? reg_csr_2079 : _GEN_2078; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2080 = 12'h820 == csr_addr[11:0] ? reg_csr_2080 : _GEN_2079; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2081 = 12'h821 == csr_addr[11:0] ? reg_csr_2081 : _GEN_2080; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2082 = 12'h822 == csr_addr[11:0] ? reg_csr_2082 : _GEN_2081; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2083 = 12'h823 == csr_addr[11:0] ? reg_csr_2083 : _GEN_2082; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2084 = 12'h824 == csr_addr[11:0] ? reg_csr_2084 : _GEN_2083; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2085 = 12'h825 == csr_addr[11:0] ? reg_csr_2085 : _GEN_2084; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2086 = 12'h826 == csr_addr[11:0] ? reg_csr_2086 : _GEN_2085; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2087 = 12'h827 == csr_addr[11:0] ? reg_csr_2087 : _GEN_2086; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2088 = 12'h828 == csr_addr[11:0] ? reg_csr_2088 : _GEN_2087; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2089 = 12'h829 == csr_addr[11:0] ? reg_csr_2089 : _GEN_2088; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2090 = 12'h82a == csr_addr[11:0] ? reg_csr_2090 : _GEN_2089; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2091 = 12'h82b == csr_addr[11:0] ? reg_csr_2091 : _GEN_2090; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2092 = 12'h82c == csr_addr[11:0] ? reg_csr_2092 : _GEN_2091; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2093 = 12'h82d == csr_addr[11:0] ? reg_csr_2093 : _GEN_2092; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2094 = 12'h82e == csr_addr[11:0] ? reg_csr_2094 : _GEN_2093; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2095 = 12'h82f == csr_addr[11:0] ? reg_csr_2095 : _GEN_2094; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2096 = 12'h830 == csr_addr[11:0] ? reg_csr_2096 : _GEN_2095; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2097 = 12'h831 == csr_addr[11:0] ? reg_csr_2097 : _GEN_2096; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2098 = 12'h832 == csr_addr[11:0] ? reg_csr_2098 : _GEN_2097; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2099 = 12'h833 == csr_addr[11:0] ? reg_csr_2099 : _GEN_2098; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2100 = 12'h834 == csr_addr[11:0] ? reg_csr_2100 : _GEN_2099; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2101 = 12'h835 == csr_addr[11:0] ? reg_csr_2101 : _GEN_2100; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2102 = 12'h836 == csr_addr[11:0] ? reg_csr_2102 : _GEN_2101; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2103 = 12'h837 == csr_addr[11:0] ? reg_csr_2103 : _GEN_2102; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2104 = 12'h838 == csr_addr[11:0] ? reg_csr_2104 : _GEN_2103; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2105 = 12'h839 == csr_addr[11:0] ? reg_csr_2105 : _GEN_2104; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2106 = 12'h83a == csr_addr[11:0] ? reg_csr_2106 : _GEN_2105; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2107 = 12'h83b == csr_addr[11:0] ? reg_csr_2107 : _GEN_2106; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2108 = 12'h83c == csr_addr[11:0] ? reg_csr_2108 : _GEN_2107; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2109 = 12'h83d == csr_addr[11:0] ? reg_csr_2109 : _GEN_2108; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2110 = 12'h83e == csr_addr[11:0] ? reg_csr_2110 : _GEN_2109; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2111 = 12'h83f == csr_addr[11:0] ? reg_csr_2111 : _GEN_2110; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2112 = 12'h840 == csr_addr[11:0] ? reg_csr_2112 : _GEN_2111; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2113 = 12'h841 == csr_addr[11:0] ? reg_csr_2113 : _GEN_2112; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2114 = 12'h842 == csr_addr[11:0] ? reg_csr_2114 : _GEN_2113; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2115 = 12'h843 == csr_addr[11:0] ? reg_csr_2115 : _GEN_2114; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2116 = 12'h844 == csr_addr[11:0] ? reg_csr_2116 : _GEN_2115; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2117 = 12'h845 == csr_addr[11:0] ? reg_csr_2117 : _GEN_2116; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2118 = 12'h846 == csr_addr[11:0] ? reg_csr_2118 : _GEN_2117; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2119 = 12'h847 == csr_addr[11:0] ? reg_csr_2119 : _GEN_2118; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2120 = 12'h848 == csr_addr[11:0] ? reg_csr_2120 : _GEN_2119; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2121 = 12'h849 == csr_addr[11:0] ? reg_csr_2121 : _GEN_2120; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2122 = 12'h84a == csr_addr[11:0] ? reg_csr_2122 : _GEN_2121; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2123 = 12'h84b == csr_addr[11:0] ? reg_csr_2123 : _GEN_2122; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2124 = 12'h84c == csr_addr[11:0] ? reg_csr_2124 : _GEN_2123; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2125 = 12'h84d == csr_addr[11:0] ? reg_csr_2125 : _GEN_2124; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2126 = 12'h84e == csr_addr[11:0] ? reg_csr_2126 : _GEN_2125; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2127 = 12'h84f == csr_addr[11:0] ? reg_csr_2127 : _GEN_2126; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2128 = 12'h850 == csr_addr[11:0] ? reg_csr_2128 : _GEN_2127; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2129 = 12'h851 == csr_addr[11:0] ? reg_csr_2129 : _GEN_2128; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2130 = 12'h852 == csr_addr[11:0] ? reg_csr_2130 : _GEN_2129; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2131 = 12'h853 == csr_addr[11:0] ? reg_csr_2131 : _GEN_2130; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2132 = 12'h854 == csr_addr[11:0] ? reg_csr_2132 : _GEN_2131; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2133 = 12'h855 == csr_addr[11:0] ? reg_csr_2133 : _GEN_2132; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2134 = 12'h856 == csr_addr[11:0] ? reg_csr_2134 : _GEN_2133; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2135 = 12'h857 == csr_addr[11:0] ? reg_csr_2135 : _GEN_2134; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2136 = 12'h858 == csr_addr[11:0] ? reg_csr_2136 : _GEN_2135; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2137 = 12'h859 == csr_addr[11:0] ? reg_csr_2137 : _GEN_2136; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2138 = 12'h85a == csr_addr[11:0] ? reg_csr_2138 : _GEN_2137; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2139 = 12'h85b == csr_addr[11:0] ? reg_csr_2139 : _GEN_2138; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2140 = 12'h85c == csr_addr[11:0] ? reg_csr_2140 : _GEN_2139; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2141 = 12'h85d == csr_addr[11:0] ? reg_csr_2141 : _GEN_2140; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2142 = 12'h85e == csr_addr[11:0] ? reg_csr_2142 : _GEN_2141; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2143 = 12'h85f == csr_addr[11:0] ? reg_csr_2143 : _GEN_2142; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2144 = 12'h860 == csr_addr[11:0] ? reg_csr_2144 : _GEN_2143; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2145 = 12'h861 == csr_addr[11:0] ? reg_csr_2145 : _GEN_2144; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2146 = 12'h862 == csr_addr[11:0] ? reg_csr_2146 : _GEN_2145; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2147 = 12'h863 == csr_addr[11:0] ? reg_csr_2147 : _GEN_2146; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2148 = 12'h864 == csr_addr[11:0] ? reg_csr_2148 : _GEN_2147; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2149 = 12'h865 == csr_addr[11:0] ? reg_csr_2149 : _GEN_2148; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2150 = 12'h866 == csr_addr[11:0] ? reg_csr_2150 : _GEN_2149; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2151 = 12'h867 == csr_addr[11:0] ? reg_csr_2151 : _GEN_2150; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2152 = 12'h868 == csr_addr[11:0] ? reg_csr_2152 : _GEN_2151; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2153 = 12'h869 == csr_addr[11:0] ? reg_csr_2153 : _GEN_2152; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2154 = 12'h86a == csr_addr[11:0] ? reg_csr_2154 : _GEN_2153; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2155 = 12'h86b == csr_addr[11:0] ? reg_csr_2155 : _GEN_2154; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2156 = 12'h86c == csr_addr[11:0] ? reg_csr_2156 : _GEN_2155; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2157 = 12'h86d == csr_addr[11:0] ? reg_csr_2157 : _GEN_2156; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2158 = 12'h86e == csr_addr[11:0] ? reg_csr_2158 : _GEN_2157; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2159 = 12'h86f == csr_addr[11:0] ? reg_csr_2159 : _GEN_2158; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2160 = 12'h870 == csr_addr[11:0] ? reg_csr_2160 : _GEN_2159; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2161 = 12'h871 == csr_addr[11:0] ? reg_csr_2161 : _GEN_2160; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2162 = 12'h872 == csr_addr[11:0] ? reg_csr_2162 : _GEN_2161; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2163 = 12'h873 == csr_addr[11:0] ? reg_csr_2163 : _GEN_2162; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2164 = 12'h874 == csr_addr[11:0] ? reg_csr_2164 : _GEN_2163; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2165 = 12'h875 == csr_addr[11:0] ? reg_csr_2165 : _GEN_2164; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2166 = 12'h876 == csr_addr[11:0] ? reg_csr_2166 : _GEN_2165; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2167 = 12'h877 == csr_addr[11:0] ? reg_csr_2167 : _GEN_2166; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2168 = 12'h878 == csr_addr[11:0] ? reg_csr_2168 : _GEN_2167; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2169 = 12'h879 == csr_addr[11:0] ? reg_csr_2169 : _GEN_2168; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2170 = 12'h87a == csr_addr[11:0] ? reg_csr_2170 : _GEN_2169; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2171 = 12'h87b == csr_addr[11:0] ? reg_csr_2171 : _GEN_2170; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2172 = 12'h87c == csr_addr[11:0] ? reg_csr_2172 : _GEN_2171; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2173 = 12'h87d == csr_addr[11:0] ? reg_csr_2173 : _GEN_2172; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2174 = 12'h87e == csr_addr[11:0] ? reg_csr_2174 : _GEN_2173; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2175 = 12'h87f == csr_addr[11:0] ? reg_csr_2175 : _GEN_2174; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2176 = 12'h880 == csr_addr[11:0] ? reg_csr_2176 : _GEN_2175; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2177 = 12'h881 == csr_addr[11:0] ? reg_csr_2177 : _GEN_2176; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2178 = 12'h882 == csr_addr[11:0] ? reg_csr_2178 : _GEN_2177; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2179 = 12'h883 == csr_addr[11:0] ? reg_csr_2179 : _GEN_2178; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2180 = 12'h884 == csr_addr[11:0] ? reg_csr_2180 : _GEN_2179; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2181 = 12'h885 == csr_addr[11:0] ? reg_csr_2181 : _GEN_2180; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2182 = 12'h886 == csr_addr[11:0] ? reg_csr_2182 : _GEN_2181; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2183 = 12'h887 == csr_addr[11:0] ? reg_csr_2183 : _GEN_2182; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2184 = 12'h888 == csr_addr[11:0] ? reg_csr_2184 : _GEN_2183; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2185 = 12'h889 == csr_addr[11:0] ? reg_csr_2185 : _GEN_2184; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2186 = 12'h88a == csr_addr[11:0] ? reg_csr_2186 : _GEN_2185; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2187 = 12'h88b == csr_addr[11:0] ? reg_csr_2187 : _GEN_2186; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2188 = 12'h88c == csr_addr[11:0] ? reg_csr_2188 : _GEN_2187; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2189 = 12'h88d == csr_addr[11:0] ? reg_csr_2189 : _GEN_2188; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2190 = 12'h88e == csr_addr[11:0] ? reg_csr_2190 : _GEN_2189; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2191 = 12'h88f == csr_addr[11:0] ? reg_csr_2191 : _GEN_2190; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2192 = 12'h890 == csr_addr[11:0] ? reg_csr_2192 : _GEN_2191; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2193 = 12'h891 == csr_addr[11:0] ? reg_csr_2193 : _GEN_2192; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2194 = 12'h892 == csr_addr[11:0] ? reg_csr_2194 : _GEN_2193; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2195 = 12'h893 == csr_addr[11:0] ? reg_csr_2195 : _GEN_2194; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2196 = 12'h894 == csr_addr[11:0] ? reg_csr_2196 : _GEN_2195; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2197 = 12'h895 == csr_addr[11:0] ? reg_csr_2197 : _GEN_2196; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2198 = 12'h896 == csr_addr[11:0] ? reg_csr_2198 : _GEN_2197; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2199 = 12'h897 == csr_addr[11:0] ? reg_csr_2199 : _GEN_2198; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2200 = 12'h898 == csr_addr[11:0] ? reg_csr_2200 : _GEN_2199; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2201 = 12'h899 == csr_addr[11:0] ? reg_csr_2201 : _GEN_2200; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2202 = 12'h89a == csr_addr[11:0] ? reg_csr_2202 : _GEN_2201; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2203 = 12'h89b == csr_addr[11:0] ? reg_csr_2203 : _GEN_2202; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2204 = 12'h89c == csr_addr[11:0] ? reg_csr_2204 : _GEN_2203; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2205 = 12'h89d == csr_addr[11:0] ? reg_csr_2205 : _GEN_2204; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2206 = 12'h89e == csr_addr[11:0] ? reg_csr_2206 : _GEN_2205; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2207 = 12'h89f == csr_addr[11:0] ? reg_csr_2207 : _GEN_2206; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2208 = 12'h8a0 == csr_addr[11:0] ? reg_csr_2208 : _GEN_2207; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2209 = 12'h8a1 == csr_addr[11:0] ? reg_csr_2209 : _GEN_2208; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2210 = 12'h8a2 == csr_addr[11:0] ? reg_csr_2210 : _GEN_2209; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2211 = 12'h8a3 == csr_addr[11:0] ? reg_csr_2211 : _GEN_2210; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2212 = 12'h8a4 == csr_addr[11:0] ? reg_csr_2212 : _GEN_2211; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2213 = 12'h8a5 == csr_addr[11:0] ? reg_csr_2213 : _GEN_2212; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2214 = 12'h8a6 == csr_addr[11:0] ? reg_csr_2214 : _GEN_2213; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2215 = 12'h8a7 == csr_addr[11:0] ? reg_csr_2215 : _GEN_2214; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2216 = 12'h8a8 == csr_addr[11:0] ? reg_csr_2216 : _GEN_2215; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2217 = 12'h8a9 == csr_addr[11:0] ? reg_csr_2217 : _GEN_2216; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2218 = 12'h8aa == csr_addr[11:0] ? reg_csr_2218 : _GEN_2217; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2219 = 12'h8ab == csr_addr[11:0] ? reg_csr_2219 : _GEN_2218; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2220 = 12'h8ac == csr_addr[11:0] ? reg_csr_2220 : _GEN_2219; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2221 = 12'h8ad == csr_addr[11:0] ? reg_csr_2221 : _GEN_2220; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2222 = 12'h8ae == csr_addr[11:0] ? reg_csr_2222 : _GEN_2221; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2223 = 12'h8af == csr_addr[11:0] ? reg_csr_2223 : _GEN_2222; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2224 = 12'h8b0 == csr_addr[11:0] ? reg_csr_2224 : _GEN_2223; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2225 = 12'h8b1 == csr_addr[11:0] ? reg_csr_2225 : _GEN_2224; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2226 = 12'h8b2 == csr_addr[11:0] ? reg_csr_2226 : _GEN_2225; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2227 = 12'h8b3 == csr_addr[11:0] ? reg_csr_2227 : _GEN_2226; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2228 = 12'h8b4 == csr_addr[11:0] ? reg_csr_2228 : _GEN_2227; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2229 = 12'h8b5 == csr_addr[11:0] ? reg_csr_2229 : _GEN_2228; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2230 = 12'h8b6 == csr_addr[11:0] ? reg_csr_2230 : _GEN_2229; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2231 = 12'h8b7 == csr_addr[11:0] ? reg_csr_2231 : _GEN_2230; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2232 = 12'h8b8 == csr_addr[11:0] ? reg_csr_2232 : _GEN_2231; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2233 = 12'h8b9 == csr_addr[11:0] ? reg_csr_2233 : _GEN_2232; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2234 = 12'h8ba == csr_addr[11:0] ? reg_csr_2234 : _GEN_2233; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2235 = 12'h8bb == csr_addr[11:0] ? reg_csr_2235 : _GEN_2234; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2236 = 12'h8bc == csr_addr[11:0] ? reg_csr_2236 : _GEN_2235; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2237 = 12'h8bd == csr_addr[11:0] ? reg_csr_2237 : _GEN_2236; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2238 = 12'h8be == csr_addr[11:0] ? reg_csr_2238 : _GEN_2237; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2239 = 12'h8bf == csr_addr[11:0] ? reg_csr_2239 : _GEN_2238; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2240 = 12'h8c0 == csr_addr[11:0] ? reg_csr_2240 : _GEN_2239; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2241 = 12'h8c1 == csr_addr[11:0] ? reg_csr_2241 : _GEN_2240; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2242 = 12'h8c2 == csr_addr[11:0] ? reg_csr_2242 : _GEN_2241; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2243 = 12'h8c3 == csr_addr[11:0] ? reg_csr_2243 : _GEN_2242; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2244 = 12'h8c4 == csr_addr[11:0] ? reg_csr_2244 : _GEN_2243; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2245 = 12'h8c5 == csr_addr[11:0] ? reg_csr_2245 : _GEN_2244; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2246 = 12'h8c6 == csr_addr[11:0] ? reg_csr_2246 : _GEN_2245; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2247 = 12'h8c7 == csr_addr[11:0] ? reg_csr_2247 : _GEN_2246; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2248 = 12'h8c8 == csr_addr[11:0] ? reg_csr_2248 : _GEN_2247; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2249 = 12'h8c9 == csr_addr[11:0] ? reg_csr_2249 : _GEN_2248; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2250 = 12'h8ca == csr_addr[11:0] ? reg_csr_2250 : _GEN_2249; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2251 = 12'h8cb == csr_addr[11:0] ? reg_csr_2251 : _GEN_2250; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2252 = 12'h8cc == csr_addr[11:0] ? reg_csr_2252 : _GEN_2251; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2253 = 12'h8cd == csr_addr[11:0] ? reg_csr_2253 : _GEN_2252; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2254 = 12'h8ce == csr_addr[11:0] ? reg_csr_2254 : _GEN_2253; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2255 = 12'h8cf == csr_addr[11:0] ? reg_csr_2255 : _GEN_2254; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2256 = 12'h8d0 == csr_addr[11:0] ? reg_csr_2256 : _GEN_2255; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2257 = 12'h8d1 == csr_addr[11:0] ? reg_csr_2257 : _GEN_2256; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2258 = 12'h8d2 == csr_addr[11:0] ? reg_csr_2258 : _GEN_2257; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2259 = 12'h8d3 == csr_addr[11:0] ? reg_csr_2259 : _GEN_2258; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2260 = 12'h8d4 == csr_addr[11:0] ? reg_csr_2260 : _GEN_2259; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2261 = 12'h8d5 == csr_addr[11:0] ? reg_csr_2261 : _GEN_2260; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2262 = 12'h8d6 == csr_addr[11:0] ? reg_csr_2262 : _GEN_2261; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2263 = 12'h8d7 == csr_addr[11:0] ? reg_csr_2263 : _GEN_2262; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2264 = 12'h8d8 == csr_addr[11:0] ? reg_csr_2264 : _GEN_2263; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2265 = 12'h8d9 == csr_addr[11:0] ? reg_csr_2265 : _GEN_2264; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2266 = 12'h8da == csr_addr[11:0] ? reg_csr_2266 : _GEN_2265; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2267 = 12'h8db == csr_addr[11:0] ? reg_csr_2267 : _GEN_2266; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2268 = 12'h8dc == csr_addr[11:0] ? reg_csr_2268 : _GEN_2267; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2269 = 12'h8dd == csr_addr[11:0] ? reg_csr_2269 : _GEN_2268; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2270 = 12'h8de == csr_addr[11:0] ? reg_csr_2270 : _GEN_2269; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2271 = 12'h8df == csr_addr[11:0] ? reg_csr_2271 : _GEN_2270; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2272 = 12'h8e0 == csr_addr[11:0] ? reg_csr_2272 : _GEN_2271; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2273 = 12'h8e1 == csr_addr[11:0] ? reg_csr_2273 : _GEN_2272; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2274 = 12'h8e2 == csr_addr[11:0] ? reg_csr_2274 : _GEN_2273; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2275 = 12'h8e3 == csr_addr[11:0] ? reg_csr_2275 : _GEN_2274; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2276 = 12'h8e4 == csr_addr[11:0] ? reg_csr_2276 : _GEN_2275; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2277 = 12'h8e5 == csr_addr[11:0] ? reg_csr_2277 : _GEN_2276; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2278 = 12'h8e6 == csr_addr[11:0] ? reg_csr_2278 : _GEN_2277; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2279 = 12'h8e7 == csr_addr[11:0] ? reg_csr_2279 : _GEN_2278; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2280 = 12'h8e8 == csr_addr[11:0] ? reg_csr_2280 : _GEN_2279; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2281 = 12'h8e9 == csr_addr[11:0] ? reg_csr_2281 : _GEN_2280; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2282 = 12'h8ea == csr_addr[11:0] ? reg_csr_2282 : _GEN_2281; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2283 = 12'h8eb == csr_addr[11:0] ? reg_csr_2283 : _GEN_2282; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2284 = 12'h8ec == csr_addr[11:0] ? reg_csr_2284 : _GEN_2283; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2285 = 12'h8ed == csr_addr[11:0] ? reg_csr_2285 : _GEN_2284; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2286 = 12'h8ee == csr_addr[11:0] ? reg_csr_2286 : _GEN_2285; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2287 = 12'h8ef == csr_addr[11:0] ? reg_csr_2287 : _GEN_2286; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2288 = 12'h8f0 == csr_addr[11:0] ? reg_csr_2288 : _GEN_2287; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2289 = 12'h8f1 == csr_addr[11:0] ? reg_csr_2289 : _GEN_2288; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2290 = 12'h8f2 == csr_addr[11:0] ? reg_csr_2290 : _GEN_2289; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2291 = 12'h8f3 == csr_addr[11:0] ? reg_csr_2291 : _GEN_2290; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2292 = 12'h8f4 == csr_addr[11:0] ? reg_csr_2292 : _GEN_2291; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2293 = 12'h8f5 == csr_addr[11:0] ? reg_csr_2293 : _GEN_2292; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2294 = 12'h8f6 == csr_addr[11:0] ? reg_csr_2294 : _GEN_2293; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2295 = 12'h8f7 == csr_addr[11:0] ? reg_csr_2295 : _GEN_2294; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2296 = 12'h8f8 == csr_addr[11:0] ? reg_csr_2296 : _GEN_2295; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2297 = 12'h8f9 == csr_addr[11:0] ? reg_csr_2297 : _GEN_2296; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2298 = 12'h8fa == csr_addr[11:0] ? reg_csr_2298 : _GEN_2297; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2299 = 12'h8fb == csr_addr[11:0] ? reg_csr_2299 : _GEN_2298; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2300 = 12'h8fc == csr_addr[11:0] ? reg_csr_2300 : _GEN_2299; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2301 = 12'h8fd == csr_addr[11:0] ? reg_csr_2301 : _GEN_2300; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2302 = 12'h8fe == csr_addr[11:0] ? reg_csr_2302 : _GEN_2301; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2303 = 12'h8ff == csr_addr[11:0] ? reg_csr_2303 : _GEN_2302; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2304 = 12'h900 == csr_addr[11:0] ? reg_csr_2304 : _GEN_2303; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2305 = 12'h901 == csr_addr[11:0] ? reg_csr_2305 : _GEN_2304; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2306 = 12'h902 == csr_addr[11:0] ? reg_csr_2306 : _GEN_2305; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2307 = 12'h903 == csr_addr[11:0] ? reg_csr_2307 : _GEN_2306; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2308 = 12'h904 == csr_addr[11:0] ? reg_csr_2308 : _GEN_2307; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2309 = 12'h905 == csr_addr[11:0] ? reg_csr_2309 : _GEN_2308; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2310 = 12'h906 == csr_addr[11:0] ? reg_csr_2310 : _GEN_2309; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2311 = 12'h907 == csr_addr[11:0] ? reg_csr_2311 : _GEN_2310; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2312 = 12'h908 == csr_addr[11:0] ? reg_csr_2312 : _GEN_2311; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2313 = 12'h909 == csr_addr[11:0] ? reg_csr_2313 : _GEN_2312; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2314 = 12'h90a == csr_addr[11:0] ? reg_csr_2314 : _GEN_2313; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2315 = 12'h90b == csr_addr[11:0] ? reg_csr_2315 : _GEN_2314; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2316 = 12'h90c == csr_addr[11:0] ? reg_csr_2316 : _GEN_2315; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2317 = 12'h90d == csr_addr[11:0] ? reg_csr_2317 : _GEN_2316; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2318 = 12'h90e == csr_addr[11:0] ? reg_csr_2318 : _GEN_2317; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2319 = 12'h90f == csr_addr[11:0] ? reg_csr_2319 : _GEN_2318; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2320 = 12'h910 == csr_addr[11:0] ? reg_csr_2320 : _GEN_2319; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2321 = 12'h911 == csr_addr[11:0] ? reg_csr_2321 : _GEN_2320; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2322 = 12'h912 == csr_addr[11:0] ? reg_csr_2322 : _GEN_2321; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2323 = 12'h913 == csr_addr[11:0] ? reg_csr_2323 : _GEN_2322; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2324 = 12'h914 == csr_addr[11:0] ? reg_csr_2324 : _GEN_2323; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2325 = 12'h915 == csr_addr[11:0] ? reg_csr_2325 : _GEN_2324; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2326 = 12'h916 == csr_addr[11:0] ? reg_csr_2326 : _GEN_2325; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2327 = 12'h917 == csr_addr[11:0] ? reg_csr_2327 : _GEN_2326; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2328 = 12'h918 == csr_addr[11:0] ? reg_csr_2328 : _GEN_2327; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2329 = 12'h919 == csr_addr[11:0] ? reg_csr_2329 : _GEN_2328; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2330 = 12'h91a == csr_addr[11:0] ? reg_csr_2330 : _GEN_2329; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2331 = 12'h91b == csr_addr[11:0] ? reg_csr_2331 : _GEN_2330; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2332 = 12'h91c == csr_addr[11:0] ? reg_csr_2332 : _GEN_2331; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2333 = 12'h91d == csr_addr[11:0] ? reg_csr_2333 : _GEN_2332; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2334 = 12'h91e == csr_addr[11:0] ? reg_csr_2334 : _GEN_2333; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2335 = 12'h91f == csr_addr[11:0] ? reg_csr_2335 : _GEN_2334; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2336 = 12'h920 == csr_addr[11:0] ? reg_csr_2336 : _GEN_2335; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2337 = 12'h921 == csr_addr[11:0] ? reg_csr_2337 : _GEN_2336; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2338 = 12'h922 == csr_addr[11:0] ? reg_csr_2338 : _GEN_2337; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2339 = 12'h923 == csr_addr[11:0] ? reg_csr_2339 : _GEN_2338; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2340 = 12'h924 == csr_addr[11:0] ? reg_csr_2340 : _GEN_2339; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2341 = 12'h925 == csr_addr[11:0] ? reg_csr_2341 : _GEN_2340; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2342 = 12'h926 == csr_addr[11:0] ? reg_csr_2342 : _GEN_2341; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2343 = 12'h927 == csr_addr[11:0] ? reg_csr_2343 : _GEN_2342; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2344 = 12'h928 == csr_addr[11:0] ? reg_csr_2344 : _GEN_2343; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2345 = 12'h929 == csr_addr[11:0] ? reg_csr_2345 : _GEN_2344; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2346 = 12'h92a == csr_addr[11:0] ? reg_csr_2346 : _GEN_2345; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2347 = 12'h92b == csr_addr[11:0] ? reg_csr_2347 : _GEN_2346; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2348 = 12'h92c == csr_addr[11:0] ? reg_csr_2348 : _GEN_2347; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2349 = 12'h92d == csr_addr[11:0] ? reg_csr_2349 : _GEN_2348; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2350 = 12'h92e == csr_addr[11:0] ? reg_csr_2350 : _GEN_2349; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2351 = 12'h92f == csr_addr[11:0] ? reg_csr_2351 : _GEN_2350; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2352 = 12'h930 == csr_addr[11:0] ? reg_csr_2352 : _GEN_2351; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2353 = 12'h931 == csr_addr[11:0] ? reg_csr_2353 : _GEN_2352; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2354 = 12'h932 == csr_addr[11:0] ? reg_csr_2354 : _GEN_2353; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2355 = 12'h933 == csr_addr[11:0] ? reg_csr_2355 : _GEN_2354; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2356 = 12'h934 == csr_addr[11:0] ? reg_csr_2356 : _GEN_2355; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2357 = 12'h935 == csr_addr[11:0] ? reg_csr_2357 : _GEN_2356; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2358 = 12'h936 == csr_addr[11:0] ? reg_csr_2358 : _GEN_2357; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2359 = 12'h937 == csr_addr[11:0] ? reg_csr_2359 : _GEN_2358; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2360 = 12'h938 == csr_addr[11:0] ? reg_csr_2360 : _GEN_2359; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2361 = 12'h939 == csr_addr[11:0] ? reg_csr_2361 : _GEN_2360; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2362 = 12'h93a == csr_addr[11:0] ? reg_csr_2362 : _GEN_2361; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2363 = 12'h93b == csr_addr[11:0] ? reg_csr_2363 : _GEN_2362; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2364 = 12'h93c == csr_addr[11:0] ? reg_csr_2364 : _GEN_2363; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2365 = 12'h93d == csr_addr[11:0] ? reg_csr_2365 : _GEN_2364; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2366 = 12'h93e == csr_addr[11:0] ? reg_csr_2366 : _GEN_2365; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2367 = 12'h93f == csr_addr[11:0] ? reg_csr_2367 : _GEN_2366; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2368 = 12'h940 == csr_addr[11:0] ? reg_csr_2368 : _GEN_2367; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2369 = 12'h941 == csr_addr[11:0] ? reg_csr_2369 : _GEN_2368; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2370 = 12'h942 == csr_addr[11:0] ? reg_csr_2370 : _GEN_2369; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2371 = 12'h943 == csr_addr[11:0] ? reg_csr_2371 : _GEN_2370; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2372 = 12'h944 == csr_addr[11:0] ? reg_csr_2372 : _GEN_2371; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2373 = 12'h945 == csr_addr[11:0] ? reg_csr_2373 : _GEN_2372; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2374 = 12'h946 == csr_addr[11:0] ? reg_csr_2374 : _GEN_2373; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2375 = 12'h947 == csr_addr[11:0] ? reg_csr_2375 : _GEN_2374; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2376 = 12'h948 == csr_addr[11:0] ? reg_csr_2376 : _GEN_2375; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2377 = 12'h949 == csr_addr[11:0] ? reg_csr_2377 : _GEN_2376; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2378 = 12'h94a == csr_addr[11:0] ? reg_csr_2378 : _GEN_2377; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2379 = 12'h94b == csr_addr[11:0] ? reg_csr_2379 : _GEN_2378; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2380 = 12'h94c == csr_addr[11:0] ? reg_csr_2380 : _GEN_2379; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2381 = 12'h94d == csr_addr[11:0] ? reg_csr_2381 : _GEN_2380; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2382 = 12'h94e == csr_addr[11:0] ? reg_csr_2382 : _GEN_2381; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2383 = 12'h94f == csr_addr[11:0] ? reg_csr_2383 : _GEN_2382; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2384 = 12'h950 == csr_addr[11:0] ? reg_csr_2384 : _GEN_2383; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2385 = 12'h951 == csr_addr[11:0] ? reg_csr_2385 : _GEN_2384; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2386 = 12'h952 == csr_addr[11:0] ? reg_csr_2386 : _GEN_2385; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2387 = 12'h953 == csr_addr[11:0] ? reg_csr_2387 : _GEN_2386; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2388 = 12'h954 == csr_addr[11:0] ? reg_csr_2388 : _GEN_2387; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2389 = 12'h955 == csr_addr[11:0] ? reg_csr_2389 : _GEN_2388; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2390 = 12'h956 == csr_addr[11:0] ? reg_csr_2390 : _GEN_2389; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2391 = 12'h957 == csr_addr[11:0] ? reg_csr_2391 : _GEN_2390; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2392 = 12'h958 == csr_addr[11:0] ? reg_csr_2392 : _GEN_2391; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2393 = 12'h959 == csr_addr[11:0] ? reg_csr_2393 : _GEN_2392; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2394 = 12'h95a == csr_addr[11:0] ? reg_csr_2394 : _GEN_2393; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2395 = 12'h95b == csr_addr[11:0] ? reg_csr_2395 : _GEN_2394; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2396 = 12'h95c == csr_addr[11:0] ? reg_csr_2396 : _GEN_2395; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2397 = 12'h95d == csr_addr[11:0] ? reg_csr_2397 : _GEN_2396; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2398 = 12'h95e == csr_addr[11:0] ? reg_csr_2398 : _GEN_2397; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2399 = 12'h95f == csr_addr[11:0] ? reg_csr_2399 : _GEN_2398; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2400 = 12'h960 == csr_addr[11:0] ? reg_csr_2400 : _GEN_2399; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2401 = 12'h961 == csr_addr[11:0] ? reg_csr_2401 : _GEN_2400; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2402 = 12'h962 == csr_addr[11:0] ? reg_csr_2402 : _GEN_2401; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2403 = 12'h963 == csr_addr[11:0] ? reg_csr_2403 : _GEN_2402; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2404 = 12'h964 == csr_addr[11:0] ? reg_csr_2404 : _GEN_2403; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2405 = 12'h965 == csr_addr[11:0] ? reg_csr_2405 : _GEN_2404; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2406 = 12'h966 == csr_addr[11:0] ? reg_csr_2406 : _GEN_2405; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2407 = 12'h967 == csr_addr[11:0] ? reg_csr_2407 : _GEN_2406; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2408 = 12'h968 == csr_addr[11:0] ? reg_csr_2408 : _GEN_2407; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2409 = 12'h969 == csr_addr[11:0] ? reg_csr_2409 : _GEN_2408; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2410 = 12'h96a == csr_addr[11:0] ? reg_csr_2410 : _GEN_2409; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2411 = 12'h96b == csr_addr[11:0] ? reg_csr_2411 : _GEN_2410; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2412 = 12'h96c == csr_addr[11:0] ? reg_csr_2412 : _GEN_2411; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2413 = 12'h96d == csr_addr[11:0] ? reg_csr_2413 : _GEN_2412; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2414 = 12'h96e == csr_addr[11:0] ? reg_csr_2414 : _GEN_2413; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2415 = 12'h96f == csr_addr[11:0] ? reg_csr_2415 : _GEN_2414; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2416 = 12'h970 == csr_addr[11:0] ? reg_csr_2416 : _GEN_2415; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2417 = 12'h971 == csr_addr[11:0] ? reg_csr_2417 : _GEN_2416; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2418 = 12'h972 == csr_addr[11:0] ? reg_csr_2418 : _GEN_2417; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2419 = 12'h973 == csr_addr[11:0] ? reg_csr_2419 : _GEN_2418; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2420 = 12'h974 == csr_addr[11:0] ? reg_csr_2420 : _GEN_2419; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2421 = 12'h975 == csr_addr[11:0] ? reg_csr_2421 : _GEN_2420; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2422 = 12'h976 == csr_addr[11:0] ? reg_csr_2422 : _GEN_2421; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2423 = 12'h977 == csr_addr[11:0] ? reg_csr_2423 : _GEN_2422; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2424 = 12'h978 == csr_addr[11:0] ? reg_csr_2424 : _GEN_2423; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2425 = 12'h979 == csr_addr[11:0] ? reg_csr_2425 : _GEN_2424; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2426 = 12'h97a == csr_addr[11:0] ? reg_csr_2426 : _GEN_2425; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2427 = 12'h97b == csr_addr[11:0] ? reg_csr_2427 : _GEN_2426; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2428 = 12'h97c == csr_addr[11:0] ? reg_csr_2428 : _GEN_2427; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2429 = 12'h97d == csr_addr[11:0] ? reg_csr_2429 : _GEN_2428; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2430 = 12'h97e == csr_addr[11:0] ? reg_csr_2430 : _GEN_2429; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2431 = 12'h97f == csr_addr[11:0] ? reg_csr_2431 : _GEN_2430; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2432 = 12'h980 == csr_addr[11:0] ? reg_csr_2432 : _GEN_2431; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2433 = 12'h981 == csr_addr[11:0] ? reg_csr_2433 : _GEN_2432; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2434 = 12'h982 == csr_addr[11:0] ? reg_csr_2434 : _GEN_2433; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2435 = 12'h983 == csr_addr[11:0] ? reg_csr_2435 : _GEN_2434; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2436 = 12'h984 == csr_addr[11:0] ? reg_csr_2436 : _GEN_2435; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2437 = 12'h985 == csr_addr[11:0] ? reg_csr_2437 : _GEN_2436; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2438 = 12'h986 == csr_addr[11:0] ? reg_csr_2438 : _GEN_2437; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2439 = 12'h987 == csr_addr[11:0] ? reg_csr_2439 : _GEN_2438; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2440 = 12'h988 == csr_addr[11:0] ? reg_csr_2440 : _GEN_2439; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2441 = 12'h989 == csr_addr[11:0] ? reg_csr_2441 : _GEN_2440; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2442 = 12'h98a == csr_addr[11:0] ? reg_csr_2442 : _GEN_2441; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2443 = 12'h98b == csr_addr[11:0] ? reg_csr_2443 : _GEN_2442; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2444 = 12'h98c == csr_addr[11:0] ? reg_csr_2444 : _GEN_2443; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2445 = 12'h98d == csr_addr[11:0] ? reg_csr_2445 : _GEN_2444; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2446 = 12'h98e == csr_addr[11:0] ? reg_csr_2446 : _GEN_2445; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2447 = 12'h98f == csr_addr[11:0] ? reg_csr_2447 : _GEN_2446; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2448 = 12'h990 == csr_addr[11:0] ? reg_csr_2448 : _GEN_2447; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2449 = 12'h991 == csr_addr[11:0] ? reg_csr_2449 : _GEN_2448; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2450 = 12'h992 == csr_addr[11:0] ? reg_csr_2450 : _GEN_2449; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2451 = 12'h993 == csr_addr[11:0] ? reg_csr_2451 : _GEN_2450; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2452 = 12'h994 == csr_addr[11:0] ? reg_csr_2452 : _GEN_2451; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2453 = 12'h995 == csr_addr[11:0] ? reg_csr_2453 : _GEN_2452; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2454 = 12'h996 == csr_addr[11:0] ? reg_csr_2454 : _GEN_2453; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2455 = 12'h997 == csr_addr[11:0] ? reg_csr_2455 : _GEN_2454; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2456 = 12'h998 == csr_addr[11:0] ? reg_csr_2456 : _GEN_2455; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2457 = 12'h999 == csr_addr[11:0] ? reg_csr_2457 : _GEN_2456; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2458 = 12'h99a == csr_addr[11:0] ? reg_csr_2458 : _GEN_2457; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2459 = 12'h99b == csr_addr[11:0] ? reg_csr_2459 : _GEN_2458; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2460 = 12'h99c == csr_addr[11:0] ? reg_csr_2460 : _GEN_2459; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2461 = 12'h99d == csr_addr[11:0] ? reg_csr_2461 : _GEN_2460; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2462 = 12'h99e == csr_addr[11:0] ? reg_csr_2462 : _GEN_2461; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2463 = 12'h99f == csr_addr[11:0] ? reg_csr_2463 : _GEN_2462; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2464 = 12'h9a0 == csr_addr[11:0] ? reg_csr_2464 : _GEN_2463; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2465 = 12'h9a1 == csr_addr[11:0] ? reg_csr_2465 : _GEN_2464; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2466 = 12'h9a2 == csr_addr[11:0] ? reg_csr_2466 : _GEN_2465; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2467 = 12'h9a3 == csr_addr[11:0] ? reg_csr_2467 : _GEN_2466; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2468 = 12'h9a4 == csr_addr[11:0] ? reg_csr_2468 : _GEN_2467; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2469 = 12'h9a5 == csr_addr[11:0] ? reg_csr_2469 : _GEN_2468; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2470 = 12'h9a6 == csr_addr[11:0] ? reg_csr_2470 : _GEN_2469; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2471 = 12'h9a7 == csr_addr[11:0] ? reg_csr_2471 : _GEN_2470; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2472 = 12'h9a8 == csr_addr[11:0] ? reg_csr_2472 : _GEN_2471; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2473 = 12'h9a9 == csr_addr[11:0] ? reg_csr_2473 : _GEN_2472; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2474 = 12'h9aa == csr_addr[11:0] ? reg_csr_2474 : _GEN_2473; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2475 = 12'h9ab == csr_addr[11:0] ? reg_csr_2475 : _GEN_2474; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2476 = 12'h9ac == csr_addr[11:0] ? reg_csr_2476 : _GEN_2475; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2477 = 12'h9ad == csr_addr[11:0] ? reg_csr_2477 : _GEN_2476; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2478 = 12'h9ae == csr_addr[11:0] ? reg_csr_2478 : _GEN_2477; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2479 = 12'h9af == csr_addr[11:0] ? reg_csr_2479 : _GEN_2478; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2480 = 12'h9b0 == csr_addr[11:0] ? reg_csr_2480 : _GEN_2479; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2481 = 12'h9b1 == csr_addr[11:0] ? reg_csr_2481 : _GEN_2480; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2482 = 12'h9b2 == csr_addr[11:0] ? reg_csr_2482 : _GEN_2481; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2483 = 12'h9b3 == csr_addr[11:0] ? reg_csr_2483 : _GEN_2482; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2484 = 12'h9b4 == csr_addr[11:0] ? reg_csr_2484 : _GEN_2483; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2485 = 12'h9b5 == csr_addr[11:0] ? reg_csr_2485 : _GEN_2484; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2486 = 12'h9b6 == csr_addr[11:0] ? reg_csr_2486 : _GEN_2485; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2487 = 12'h9b7 == csr_addr[11:0] ? reg_csr_2487 : _GEN_2486; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2488 = 12'h9b8 == csr_addr[11:0] ? reg_csr_2488 : _GEN_2487; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2489 = 12'h9b9 == csr_addr[11:0] ? reg_csr_2489 : _GEN_2488; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2490 = 12'h9ba == csr_addr[11:0] ? reg_csr_2490 : _GEN_2489; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2491 = 12'h9bb == csr_addr[11:0] ? reg_csr_2491 : _GEN_2490; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2492 = 12'h9bc == csr_addr[11:0] ? reg_csr_2492 : _GEN_2491; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2493 = 12'h9bd == csr_addr[11:0] ? reg_csr_2493 : _GEN_2492; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2494 = 12'h9be == csr_addr[11:0] ? reg_csr_2494 : _GEN_2493; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2495 = 12'h9bf == csr_addr[11:0] ? reg_csr_2495 : _GEN_2494; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2496 = 12'h9c0 == csr_addr[11:0] ? reg_csr_2496 : _GEN_2495; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2497 = 12'h9c1 == csr_addr[11:0] ? reg_csr_2497 : _GEN_2496; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2498 = 12'h9c2 == csr_addr[11:0] ? reg_csr_2498 : _GEN_2497; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2499 = 12'h9c3 == csr_addr[11:0] ? reg_csr_2499 : _GEN_2498; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2500 = 12'h9c4 == csr_addr[11:0] ? reg_csr_2500 : _GEN_2499; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2501 = 12'h9c5 == csr_addr[11:0] ? reg_csr_2501 : _GEN_2500; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2502 = 12'h9c6 == csr_addr[11:0] ? reg_csr_2502 : _GEN_2501; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2503 = 12'h9c7 == csr_addr[11:0] ? reg_csr_2503 : _GEN_2502; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2504 = 12'h9c8 == csr_addr[11:0] ? reg_csr_2504 : _GEN_2503; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2505 = 12'h9c9 == csr_addr[11:0] ? reg_csr_2505 : _GEN_2504; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2506 = 12'h9ca == csr_addr[11:0] ? reg_csr_2506 : _GEN_2505; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2507 = 12'h9cb == csr_addr[11:0] ? reg_csr_2507 : _GEN_2506; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2508 = 12'h9cc == csr_addr[11:0] ? reg_csr_2508 : _GEN_2507; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2509 = 12'h9cd == csr_addr[11:0] ? reg_csr_2509 : _GEN_2508; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2510 = 12'h9ce == csr_addr[11:0] ? reg_csr_2510 : _GEN_2509; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2511 = 12'h9cf == csr_addr[11:0] ? reg_csr_2511 : _GEN_2510; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2512 = 12'h9d0 == csr_addr[11:0] ? reg_csr_2512 : _GEN_2511; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2513 = 12'h9d1 == csr_addr[11:0] ? reg_csr_2513 : _GEN_2512; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2514 = 12'h9d2 == csr_addr[11:0] ? reg_csr_2514 : _GEN_2513; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2515 = 12'h9d3 == csr_addr[11:0] ? reg_csr_2515 : _GEN_2514; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2516 = 12'h9d4 == csr_addr[11:0] ? reg_csr_2516 : _GEN_2515; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2517 = 12'h9d5 == csr_addr[11:0] ? reg_csr_2517 : _GEN_2516; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2518 = 12'h9d6 == csr_addr[11:0] ? reg_csr_2518 : _GEN_2517; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2519 = 12'h9d7 == csr_addr[11:0] ? reg_csr_2519 : _GEN_2518; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2520 = 12'h9d8 == csr_addr[11:0] ? reg_csr_2520 : _GEN_2519; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2521 = 12'h9d9 == csr_addr[11:0] ? reg_csr_2521 : _GEN_2520; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2522 = 12'h9da == csr_addr[11:0] ? reg_csr_2522 : _GEN_2521; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2523 = 12'h9db == csr_addr[11:0] ? reg_csr_2523 : _GEN_2522; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2524 = 12'h9dc == csr_addr[11:0] ? reg_csr_2524 : _GEN_2523; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2525 = 12'h9dd == csr_addr[11:0] ? reg_csr_2525 : _GEN_2524; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2526 = 12'h9de == csr_addr[11:0] ? reg_csr_2526 : _GEN_2525; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2527 = 12'h9df == csr_addr[11:0] ? reg_csr_2527 : _GEN_2526; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2528 = 12'h9e0 == csr_addr[11:0] ? reg_csr_2528 : _GEN_2527; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2529 = 12'h9e1 == csr_addr[11:0] ? reg_csr_2529 : _GEN_2528; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2530 = 12'h9e2 == csr_addr[11:0] ? reg_csr_2530 : _GEN_2529; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2531 = 12'h9e3 == csr_addr[11:0] ? reg_csr_2531 : _GEN_2530; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2532 = 12'h9e4 == csr_addr[11:0] ? reg_csr_2532 : _GEN_2531; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2533 = 12'h9e5 == csr_addr[11:0] ? reg_csr_2533 : _GEN_2532; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2534 = 12'h9e6 == csr_addr[11:0] ? reg_csr_2534 : _GEN_2533; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2535 = 12'h9e7 == csr_addr[11:0] ? reg_csr_2535 : _GEN_2534; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2536 = 12'h9e8 == csr_addr[11:0] ? reg_csr_2536 : _GEN_2535; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2537 = 12'h9e9 == csr_addr[11:0] ? reg_csr_2537 : _GEN_2536; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2538 = 12'h9ea == csr_addr[11:0] ? reg_csr_2538 : _GEN_2537; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2539 = 12'h9eb == csr_addr[11:0] ? reg_csr_2539 : _GEN_2538; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2540 = 12'h9ec == csr_addr[11:0] ? reg_csr_2540 : _GEN_2539; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2541 = 12'h9ed == csr_addr[11:0] ? reg_csr_2541 : _GEN_2540; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2542 = 12'h9ee == csr_addr[11:0] ? reg_csr_2542 : _GEN_2541; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2543 = 12'h9ef == csr_addr[11:0] ? reg_csr_2543 : _GEN_2542; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2544 = 12'h9f0 == csr_addr[11:0] ? reg_csr_2544 : _GEN_2543; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2545 = 12'h9f1 == csr_addr[11:0] ? reg_csr_2545 : _GEN_2544; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2546 = 12'h9f2 == csr_addr[11:0] ? reg_csr_2546 : _GEN_2545; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2547 = 12'h9f3 == csr_addr[11:0] ? reg_csr_2547 : _GEN_2546; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2548 = 12'h9f4 == csr_addr[11:0] ? reg_csr_2548 : _GEN_2547; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2549 = 12'h9f5 == csr_addr[11:0] ? reg_csr_2549 : _GEN_2548; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2550 = 12'h9f6 == csr_addr[11:0] ? reg_csr_2550 : _GEN_2549; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2551 = 12'h9f7 == csr_addr[11:0] ? reg_csr_2551 : _GEN_2550; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2552 = 12'h9f8 == csr_addr[11:0] ? reg_csr_2552 : _GEN_2551; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2553 = 12'h9f9 == csr_addr[11:0] ? reg_csr_2553 : _GEN_2552; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2554 = 12'h9fa == csr_addr[11:0] ? reg_csr_2554 : _GEN_2553; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2555 = 12'h9fb == csr_addr[11:0] ? reg_csr_2555 : _GEN_2554; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2556 = 12'h9fc == csr_addr[11:0] ? reg_csr_2556 : _GEN_2555; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2557 = 12'h9fd == csr_addr[11:0] ? reg_csr_2557 : _GEN_2556; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2558 = 12'h9fe == csr_addr[11:0] ? reg_csr_2558 : _GEN_2557; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2559 = 12'h9ff == csr_addr[11:0] ? reg_csr_2559 : _GEN_2558; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2560 = 12'ha00 == csr_addr[11:0] ? reg_csr_2560 : _GEN_2559; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2561 = 12'ha01 == csr_addr[11:0] ? reg_csr_2561 : _GEN_2560; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2562 = 12'ha02 == csr_addr[11:0] ? reg_csr_2562 : _GEN_2561; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2563 = 12'ha03 == csr_addr[11:0] ? reg_csr_2563 : _GEN_2562; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2564 = 12'ha04 == csr_addr[11:0] ? reg_csr_2564 : _GEN_2563; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2565 = 12'ha05 == csr_addr[11:0] ? reg_csr_2565 : _GEN_2564; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2566 = 12'ha06 == csr_addr[11:0] ? reg_csr_2566 : _GEN_2565; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2567 = 12'ha07 == csr_addr[11:0] ? reg_csr_2567 : _GEN_2566; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2568 = 12'ha08 == csr_addr[11:0] ? reg_csr_2568 : _GEN_2567; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2569 = 12'ha09 == csr_addr[11:0] ? reg_csr_2569 : _GEN_2568; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2570 = 12'ha0a == csr_addr[11:0] ? reg_csr_2570 : _GEN_2569; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2571 = 12'ha0b == csr_addr[11:0] ? reg_csr_2571 : _GEN_2570; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2572 = 12'ha0c == csr_addr[11:0] ? reg_csr_2572 : _GEN_2571; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2573 = 12'ha0d == csr_addr[11:0] ? reg_csr_2573 : _GEN_2572; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2574 = 12'ha0e == csr_addr[11:0] ? reg_csr_2574 : _GEN_2573; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2575 = 12'ha0f == csr_addr[11:0] ? reg_csr_2575 : _GEN_2574; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2576 = 12'ha10 == csr_addr[11:0] ? reg_csr_2576 : _GEN_2575; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2577 = 12'ha11 == csr_addr[11:0] ? reg_csr_2577 : _GEN_2576; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2578 = 12'ha12 == csr_addr[11:0] ? reg_csr_2578 : _GEN_2577; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2579 = 12'ha13 == csr_addr[11:0] ? reg_csr_2579 : _GEN_2578; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2580 = 12'ha14 == csr_addr[11:0] ? reg_csr_2580 : _GEN_2579; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2581 = 12'ha15 == csr_addr[11:0] ? reg_csr_2581 : _GEN_2580; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2582 = 12'ha16 == csr_addr[11:0] ? reg_csr_2582 : _GEN_2581; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2583 = 12'ha17 == csr_addr[11:0] ? reg_csr_2583 : _GEN_2582; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2584 = 12'ha18 == csr_addr[11:0] ? reg_csr_2584 : _GEN_2583; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2585 = 12'ha19 == csr_addr[11:0] ? reg_csr_2585 : _GEN_2584; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2586 = 12'ha1a == csr_addr[11:0] ? reg_csr_2586 : _GEN_2585; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2587 = 12'ha1b == csr_addr[11:0] ? reg_csr_2587 : _GEN_2586; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2588 = 12'ha1c == csr_addr[11:0] ? reg_csr_2588 : _GEN_2587; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2589 = 12'ha1d == csr_addr[11:0] ? reg_csr_2589 : _GEN_2588; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2590 = 12'ha1e == csr_addr[11:0] ? reg_csr_2590 : _GEN_2589; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2591 = 12'ha1f == csr_addr[11:0] ? reg_csr_2591 : _GEN_2590; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2592 = 12'ha20 == csr_addr[11:0] ? reg_csr_2592 : _GEN_2591; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2593 = 12'ha21 == csr_addr[11:0] ? reg_csr_2593 : _GEN_2592; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2594 = 12'ha22 == csr_addr[11:0] ? reg_csr_2594 : _GEN_2593; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2595 = 12'ha23 == csr_addr[11:0] ? reg_csr_2595 : _GEN_2594; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2596 = 12'ha24 == csr_addr[11:0] ? reg_csr_2596 : _GEN_2595; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2597 = 12'ha25 == csr_addr[11:0] ? reg_csr_2597 : _GEN_2596; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2598 = 12'ha26 == csr_addr[11:0] ? reg_csr_2598 : _GEN_2597; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2599 = 12'ha27 == csr_addr[11:0] ? reg_csr_2599 : _GEN_2598; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2600 = 12'ha28 == csr_addr[11:0] ? reg_csr_2600 : _GEN_2599; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2601 = 12'ha29 == csr_addr[11:0] ? reg_csr_2601 : _GEN_2600; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2602 = 12'ha2a == csr_addr[11:0] ? reg_csr_2602 : _GEN_2601; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2603 = 12'ha2b == csr_addr[11:0] ? reg_csr_2603 : _GEN_2602; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2604 = 12'ha2c == csr_addr[11:0] ? reg_csr_2604 : _GEN_2603; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2605 = 12'ha2d == csr_addr[11:0] ? reg_csr_2605 : _GEN_2604; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2606 = 12'ha2e == csr_addr[11:0] ? reg_csr_2606 : _GEN_2605; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2607 = 12'ha2f == csr_addr[11:0] ? reg_csr_2607 : _GEN_2606; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2608 = 12'ha30 == csr_addr[11:0] ? reg_csr_2608 : _GEN_2607; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2609 = 12'ha31 == csr_addr[11:0] ? reg_csr_2609 : _GEN_2608; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2610 = 12'ha32 == csr_addr[11:0] ? reg_csr_2610 : _GEN_2609; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2611 = 12'ha33 == csr_addr[11:0] ? reg_csr_2611 : _GEN_2610; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2612 = 12'ha34 == csr_addr[11:0] ? reg_csr_2612 : _GEN_2611; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2613 = 12'ha35 == csr_addr[11:0] ? reg_csr_2613 : _GEN_2612; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2614 = 12'ha36 == csr_addr[11:0] ? reg_csr_2614 : _GEN_2613; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2615 = 12'ha37 == csr_addr[11:0] ? reg_csr_2615 : _GEN_2614; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2616 = 12'ha38 == csr_addr[11:0] ? reg_csr_2616 : _GEN_2615; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2617 = 12'ha39 == csr_addr[11:0] ? reg_csr_2617 : _GEN_2616; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2618 = 12'ha3a == csr_addr[11:0] ? reg_csr_2618 : _GEN_2617; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2619 = 12'ha3b == csr_addr[11:0] ? reg_csr_2619 : _GEN_2618; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2620 = 12'ha3c == csr_addr[11:0] ? reg_csr_2620 : _GEN_2619; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2621 = 12'ha3d == csr_addr[11:0] ? reg_csr_2621 : _GEN_2620; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2622 = 12'ha3e == csr_addr[11:0] ? reg_csr_2622 : _GEN_2621; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2623 = 12'ha3f == csr_addr[11:0] ? reg_csr_2623 : _GEN_2622; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2624 = 12'ha40 == csr_addr[11:0] ? reg_csr_2624 : _GEN_2623; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2625 = 12'ha41 == csr_addr[11:0] ? reg_csr_2625 : _GEN_2624; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2626 = 12'ha42 == csr_addr[11:0] ? reg_csr_2626 : _GEN_2625; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2627 = 12'ha43 == csr_addr[11:0] ? reg_csr_2627 : _GEN_2626; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2628 = 12'ha44 == csr_addr[11:0] ? reg_csr_2628 : _GEN_2627; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2629 = 12'ha45 == csr_addr[11:0] ? reg_csr_2629 : _GEN_2628; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2630 = 12'ha46 == csr_addr[11:0] ? reg_csr_2630 : _GEN_2629; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2631 = 12'ha47 == csr_addr[11:0] ? reg_csr_2631 : _GEN_2630; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2632 = 12'ha48 == csr_addr[11:0] ? reg_csr_2632 : _GEN_2631; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2633 = 12'ha49 == csr_addr[11:0] ? reg_csr_2633 : _GEN_2632; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2634 = 12'ha4a == csr_addr[11:0] ? reg_csr_2634 : _GEN_2633; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2635 = 12'ha4b == csr_addr[11:0] ? reg_csr_2635 : _GEN_2634; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2636 = 12'ha4c == csr_addr[11:0] ? reg_csr_2636 : _GEN_2635; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2637 = 12'ha4d == csr_addr[11:0] ? reg_csr_2637 : _GEN_2636; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2638 = 12'ha4e == csr_addr[11:0] ? reg_csr_2638 : _GEN_2637; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2639 = 12'ha4f == csr_addr[11:0] ? reg_csr_2639 : _GEN_2638; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2640 = 12'ha50 == csr_addr[11:0] ? reg_csr_2640 : _GEN_2639; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2641 = 12'ha51 == csr_addr[11:0] ? reg_csr_2641 : _GEN_2640; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2642 = 12'ha52 == csr_addr[11:0] ? reg_csr_2642 : _GEN_2641; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2643 = 12'ha53 == csr_addr[11:0] ? reg_csr_2643 : _GEN_2642; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2644 = 12'ha54 == csr_addr[11:0] ? reg_csr_2644 : _GEN_2643; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2645 = 12'ha55 == csr_addr[11:0] ? reg_csr_2645 : _GEN_2644; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2646 = 12'ha56 == csr_addr[11:0] ? reg_csr_2646 : _GEN_2645; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2647 = 12'ha57 == csr_addr[11:0] ? reg_csr_2647 : _GEN_2646; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2648 = 12'ha58 == csr_addr[11:0] ? reg_csr_2648 : _GEN_2647; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2649 = 12'ha59 == csr_addr[11:0] ? reg_csr_2649 : _GEN_2648; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2650 = 12'ha5a == csr_addr[11:0] ? reg_csr_2650 : _GEN_2649; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2651 = 12'ha5b == csr_addr[11:0] ? reg_csr_2651 : _GEN_2650; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2652 = 12'ha5c == csr_addr[11:0] ? reg_csr_2652 : _GEN_2651; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2653 = 12'ha5d == csr_addr[11:0] ? reg_csr_2653 : _GEN_2652; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2654 = 12'ha5e == csr_addr[11:0] ? reg_csr_2654 : _GEN_2653; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2655 = 12'ha5f == csr_addr[11:0] ? reg_csr_2655 : _GEN_2654; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2656 = 12'ha60 == csr_addr[11:0] ? reg_csr_2656 : _GEN_2655; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2657 = 12'ha61 == csr_addr[11:0] ? reg_csr_2657 : _GEN_2656; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2658 = 12'ha62 == csr_addr[11:0] ? reg_csr_2658 : _GEN_2657; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2659 = 12'ha63 == csr_addr[11:0] ? reg_csr_2659 : _GEN_2658; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2660 = 12'ha64 == csr_addr[11:0] ? reg_csr_2660 : _GEN_2659; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2661 = 12'ha65 == csr_addr[11:0] ? reg_csr_2661 : _GEN_2660; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2662 = 12'ha66 == csr_addr[11:0] ? reg_csr_2662 : _GEN_2661; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2663 = 12'ha67 == csr_addr[11:0] ? reg_csr_2663 : _GEN_2662; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2664 = 12'ha68 == csr_addr[11:0] ? reg_csr_2664 : _GEN_2663; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2665 = 12'ha69 == csr_addr[11:0] ? reg_csr_2665 : _GEN_2664; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2666 = 12'ha6a == csr_addr[11:0] ? reg_csr_2666 : _GEN_2665; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2667 = 12'ha6b == csr_addr[11:0] ? reg_csr_2667 : _GEN_2666; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2668 = 12'ha6c == csr_addr[11:0] ? reg_csr_2668 : _GEN_2667; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2669 = 12'ha6d == csr_addr[11:0] ? reg_csr_2669 : _GEN_2668; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2670 = 12'ha6e == csr_addr[11:0] ? reg_csr_2670 : _GEN_2669; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2671 = 12'ha6f == csr_addr[11:0] ? reg_csr_2671 : _GEN_2670; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2672 = 12'ha70 == csr_addr[11:0] ? reg_csr_2672 : _GEN_2671; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2673 = 12'ha71 == csr_addr[11:0] ? reg_csr_2673 : _GEN_2672; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2674 = 12'ha72 == csr_addr[11:0] ? reg_csr_2674 : _GEN_2673; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2675 = 12'ha73 == csr_addr[11:0] ? reg_csr_2675 : _GEN_2674; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2676 = 12'ha74 == csr_addr[11:0] ? reg_csr_2676 : _GEN_2675; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2677 = 12'ha75 == csr_addr[11:0] ? reg_csr_2677 : _GEN_2676; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2678 = 12'ha76 == csr_addr[11:0] ? reg_csr_2678 : _GEN_2677; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2679 = 12'ha77 == csr_addr[11:0] ? reg_csr_2679 : _GEN_2678; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2680 = 12'ha78 == csr_addr[11:0] ? reg_csr_2680 : _GEN_2679; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2681 = 12'ha79 == csr_addr[11:0] ? reg_csr_2681 : _GEN_2680; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2682 = 12'ha7a == csr_addr[11:0] ? reg_csr_2682 : _GEN_2681; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2683 = 12'ha7b == csr_addr[11:0] ? reg_csr_2683 : _GEN_2682; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2684 = 12'ha7c == csr_addr[11:0] ? reg_csr_2684 : _GEN_2683; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2685 = 12'ha7d == csr_addr[11:0] ? reg_csr_2685 : _GEN_2684; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2686 = 12'ha7e == csr_addr[11:0] ? reg_csr_2686 : _GEN_2685; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2687 = 12'ha7f == csr_addr[11:0] ? reg_csr_2687 : _GEN_2686; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2688 = 12'ha80 == csr_addr[11:0] ? reg_csr_2688 : _GEN_2687; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2689 = 12'ha81 == csr_addr[11:0] ? reg_csr_2689 : _GEN_2688; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2690 = 12'ha82 == csr_addr[11:0] ? reg_csr_2690 : _GEN_2689; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2691 = 12'ha83 == csr_addr[11:0] ? reg_csr_2691 : _GEN_2690; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2692 = 12'ha84 == csr_addr[11:0] ? reg_csr_2692 : _GEN_2691; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2693 = 12'ha85 == csr_addr[11:0] ? reg_csr_2693 : _GEN_2692; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2694 = 12'ha86 == csr_addr[11:0] ? reg_csr_2694 : _GEN_2693; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2695 = 12'ha87 == csr_addr[11:0] ? reg_csr_2695 : _GEN_2694; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2696 = 12'ha88 == csr_addr[11:0] ? reg_csr_2696 : _GEN_2695; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2697 = 12'ha89 == csr_addr[11:0] ? reg_csr_2697 : _GEN_2696; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2698 = 12'ha8a == csr_addr[11:0] ? reg_csr_2698 : _GEN_2697; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2699 = 12'ha8b == csr_addr[11:0] ? reg_csr_2699 : _GEN_2698; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2700 = 12'ha8c == csr_addr[11:0] ? reg_csr_2700 : _GEN_2699; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2701 = 12'ha8d == csr_addr[11:0] ? reg_csr_2701 : _GEN_2700; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2702 = 12'ha8e == csr_addr[11:0] ? reg_csr_2702 : _GEN_2701; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2703 = 12'ha8f == csr_addr[11:0] ? reg_csr_2703 : _GEN_2702; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2704 = 12'ha90 == csr_addr[11:0] ? reg_csr_2704 : _GEN_2703; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2705 = 12'ha91 == csr_addr[11:0] ? reg_csr_2705 : _GEN_2704; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2706 = 12'ha92 == csr_addr[11:0] ? reg_csr_2706 : _GEN_2705; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2707 = 12'ha93 == csr_addr[11:0] ? reg_csr_2707 : _GEN_2706; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2708 = 12'ha94 == csr_addr[11:0] ? reg_csr_2708 : _GEN_2707; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2709 = 12'ha95 == csr_addr[11:0] ? reg_csr_2709 : _GEN_2708; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2710 = 12'ha96 == csr_addr[11:0] ? reg_csr_2710 : _GEN_2709; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2711 = 12'ha97 == csr_addr[11:0] ? reg_csr_2711 : _GEN_2710; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2712 = 12'ha98 == csr_addr[11:0] ? reg_csr_2712 : _GEN_2711; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2713 = 12'ha99 == csr_addr[11:0] ? reg_csr_2713 : _GEN_2712; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2714 = 12'ha9a == csr_addr[11:0] ? reg_csr_2714 : _GEN_2713; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2715 = 12'ha9b == csr_addr[11:0] ? reg_csr_2715 : _GEN_2714; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2716 = 12'ha9c == csr_addr[11:0] ? reg_csr_2716 : _GEN_2715; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2717 = 12'ha9d == csr_addr[11:0] ? reg_csr_2717 : _GEN_2716; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2718 = 12'ha9e == csr_addr[11:0] ? reg_csr_2718 : _GEN_2717; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2719 = 12'ha9f == csr_addr[11:0] ? reg_csr_2719 : _GEN_2718; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2720 = 12'haa0 == csr_addr[11:0] ? reg_csr_2720 : _GEN_2719; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2721 = 12'haa1 == csr_addr[11:0] ? reg_csr_2721 : _GEN_2720; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2722 = 12'haa2 == csr_addr[11:0] ? reg_csr_2722 : _GEN_2721; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2723 = 12'haa3 == csr_addr[11:0] ? reg_csr_2723 : _GEN_2722; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2724 = 12'haa4 == csr_addr[11:0] ? reg_csr_2724 : _GEN_2723; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2725 = 12'haa5 == csr_addr[11:0] ? reg_csr_2725 : _GEN_2724; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2726 = 12'haa6 == csr_addr[11:0] ? reg_csr_2726 : _GEN_2725; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2727 = 12'haa7 == csr_addr[11:0] ? reg_csr_2727 : _GEN_2726; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2728 = 12'haa8 == csr_addr[11:0] ? reg_csr_2728 : _GEN_2727; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2729 = 12'haa9 == csr_addr[11:0] ? reg_csr_2729 : _GEN_2728; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2730 = 12'haaa == csr_addr[11:0] ? reg_csr_2730 : _GEN_2729; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2731 = 12'haab == csr_addr[11:0] ? reg_csr_2731 : _GEN_2730; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2732 = 12'haac == csr_addr[11:0] ? reg_csr_2732 : _GEN_2731; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2733 = 12'haad == csr_addr[11:0] ? reg_csr_2733 : _GEN_2732; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2734 = 12'haae == csr_addr[11:0] ? reg_csr_2734 : _GEN_2733; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2735 = 12'haaf == csr_addr[11:0] ? reg_csr_2735 : _GEN_2734; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2736 = 12'hab0 == csr_addr[11:0] ? reg_csr_2736 : _GEN_2735; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2737 = 12'hab1 == csr_addr[11:0] ? reg_csr_2737 : _GEN_2736; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2738 = 12'hab2 == csr_addr[11:0] ? reg_csr_2738 : _GEN_2737; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2739 = 12'hab3 == csr_addr[11:0] ? reg_csr_2739 : _GEN_2738; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2740 = 12'hab4 == csr_addr[11:0] ? reg_csr_2740 : _GEN_2739; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2741 = 12'hab5 == csr_addr[11:0] ? reg_csr_2741 : _GEN_2740; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2742 = 12'hab6 == csr_addr[11:0] ? reg_csr_2742 : _GEN_2741; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2743 = 12'hab7 == csr_addr[11:0] ? reg_csr_2743 : _GEN_2742; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2744 = 12'hab8 == csr_addr[11:0] ? reg_csr_2744 : _GEN_2743; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2745 = 12'hab9 == csr_addr[11:0] ? reg_csr_2745 : _GEN_2744; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2746 = 12'haba == csr_addr[11:0] ? reg_csr_2746 : _GEN_2745; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2747 = 12'habb == csr_addr[11:0] ? reg_csr_2747 : _GEN_2746; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2748 = 12'habc == csr_addr[11:0] ? reg_csr_2748 : _GEN_2747; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2749 = 12'habd == csr_addr[11:0] ? reg_csr_2749 : _GEN_2748; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2750 = 12'habe == csr_addr[11:0] ? reg_csr_2750 : _GEN_2749; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2751 = 12'habf == csr_addr[11:0] ? reg_csr_2751 : _GEN_2750; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2752 = 12'hac0 == csr_addr[11:0] ? reg_csr_2752 : _GEN_2751; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2753 = 12'hac1 == csr_addr[11:0] ? reg_csr_2753 : _GEN_2752; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2754 = 12'hac2 == csr_addr[11:0] ? reg_csr_2754 : _GEN_2753; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2755 = 12'hac3 == csr_addr[11:0] ? reg_csr_2755 : _GEN_2754; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2756 = 12'hac4 == csr_addr[11:0] ? reg_csr_2756 : _GEN_2755; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2757 = 12'hac5 == csr_addr[11:0] ? reg_csr_2757 : _GEN_2756; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2758 = 12'hac6 == csr_addr[11:0] ? reg_csr_2758 : _GEN_2757; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2759 = 12'hac7 == csr_addr[11:0] ? reg_csr_2759 : _GEN_2758; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2760 = 12'hac8 == csr_addr[11:0] ? reg_csr_2760 : _GEN_2759; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2761 = 12'hac9 == csr_addr[11:0] ? reg_csr_2761 : _GEN_2760; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2762 = 12'haca == csr_addr[11:0] ? reg_csr_2762 : _GEN_2761; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2763 = 12'hacb == csr_addr[11:0] ? reg_csr_2763 : _GEN_2762; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2764 = 12'hacc == csr_addr[11:0] ? reg_csr_2764 : _GEN_2763; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2765 = 12'hacd == csr_addr[11:0] ? reg_csr_2765 : _GEN_2764; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2766 = 12'hace == csr_addr[11:0] ? reg_csr_2766 : _GEN_2765; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2767 = 12'hacf == csr_addr[11:0] ? reg_csr_2767 : _GEN_2766; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2768 = 12'had0 == csr_addr[11:0] ? reg_csr_2768 : _GEN_2767; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2769 = 12'had1 == csr_addr[11:0] ? reg_csr_2769 : _GEN_2768; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2770 = 12'had2 == csr_addr[11:0] ? reg_csr_2770 : _GEN_2769; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2771 = 12'had3 == csr_addr[11:0] ? reg_csr_2771 : _GEN_2770; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2772 = 12'had4 == csr_addr[11:0] ? reg_csr_2772 : _GEN_2771; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2773 = 12'had5 == csr_addr[11:0] ? reg_csr_2773 : _GEN_2772; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2774 = 12'had6 == csr_addr[11:0] ? reg_csr_2774 : _GEN_2773; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2775 = 12'had7 == csr_addr[11:0] ? reg_csr_2775 : _GEN_2774; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2776 = 12'had8 == csr_addr[11:0] ? reg_csr_2776 : _GEN_2775; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2777 = 12'had9 == csr_addr[11:0] ? reg_csr_2777 : _GEN_2776; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2778 = 12'hada == csr_addr[11:0] ? reg_csr_2778 : _GEN_2777; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2779 = 12'hadb == csr_addr[11:0] ? reg_csr_2779 : _GEN_2778; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2780 = 12'hadc == csr_addr[11:0] ? reg_csr_2780 : _GEN_2779; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2781 = 12'hadd == csr_addr[11:0] ? reg_csr_2781 : _GEN_2780; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2782 = 12'hade == csr_addr[11:0] ? reg_csr_2782 : _GEN_2781; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2783 = 12'hadf == csr_addr[11:0] ? reg_csr_2783 : _GEN_2782; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2784 = 12'hae0 == csr_addr[11:0] ? reg_csr_2784 : _GEN_2783; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2785 = 12'hae1 == csr_addr[11:0] ? reg_csr_2785 : _GEN_2784; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2786 = 12'hae2 == csr_addr[11:0] ? reg_csr_2786 : _GEN_2785; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2787 = 12'hae3 == csr_addr[11:0] ? reg_csr_2787 : _GEN_2786; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2788 = 12'hae4 == csr_addr[11:0] ? reg_csr_2788 : _GEN_2787; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2789 = 12'hae5 == csr_addr[11:0] ? reg_csr_2789 : _GEN_2788; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2790 = 12'hae6 == csr_addr[11:0] ? reg_csr_2790 : _GEN_2789; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2791 = 12'hae7 == csr_addr[11:0] ? reg_csr_2791 : _GEN_2790; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2792 = 12'hae8 == csr_addr[11:0] ? reg_csr_2792 : _GEN_2791; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2793 = 12'hae9 == csr_addr[11:0] ? reg_csr_2793 : _GEN_2792; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2794 = 12'haea == csr_addr[11:0] ? reg_csr_2794 : _GEN_2793; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2795 = 12'haeb == csr_addr[11:0] ? reg_csr_2795 : _GEN_2794; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2796 = 12'haec == csr_addr[11:0] ? reg_csr_2796 : _GEN_2795; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2797 = 12'haed == csr_addr[11:0] ? reg_csr_2797 : _GEN_2796; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2798 = 12'haee == csr_addr[11:0] ? reg_csr_2798 : _GEN_2797; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2799 = 12'haef == csr_addr[11:0] ? reg_csr_2799 : _GEN_2798; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2800 = 12'haf0 == csr_addr[11:0] ? reg_csr_2800 : _GEN_2799; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2801 = 12'haf1 == csr_addr[11:0] ? reg_csr_2801 : _GEN_2800; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2802 = 12'haf2 == csr_addr[11:0] ? reg_csr_2802 : _GEN_2801; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2803 = 12'haf3 == csr_addr[11:0] ? reg_csr_2803 : _GEN_2802; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2804 = 12'haf4 == csr_addr[11:0] ? reg_csr_2804 : _GEN_2803; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2805 = 12'haf5 == csr_addr[11:0] ? reg_csr_2805 : _GEN_2804; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2806 = 12'haf6 == csr_addr[11:0] ? reg_csr_2806 : _GEN_2805; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2807 = 12'haf7 == csr_addr[11:0] ? reg_csr_2807 : _GEN_2806; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2808 = 12'haf8 == csr_addr[11:0] ? reg_csr_2808 : _GEN_2807; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2809 = 12'haf9 == csr_addr[11:0] ? reg_csr_2809 : _GEN_2808; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2810 = 12'hafa == csr_addr[11:0] ? reg_csr_2810 : _GEN_2809; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2811 = 12'hafb == csr_addr[11:0] ? reg_csr_2811 : _GEN_2810; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2812 = 12'hafc == csr_addr[11:0] ? reg_csr_2812 : _GEN_2811; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2813 = 12'hafd == csr_addr[11:0] ? reg_csr_2813 : _GEN_2812; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2814 = 12'hafe == csr_addr[11:0] ? reg_csr_2814 : _GEN_2813; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2815 = 12'haff == csr_addr[11:0] ? reg_csr_2815 : _GEN_2814; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2816 = 12'hb00 == csr_addr[11:0] ? reg_csr_2816 : _GEN_2815; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2817 = 12'hb01 == csr_addr[11:0] ? reg_csr_2817 : _GEN_2816; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2818 = 12'hb02 == csr_addr[11:0] ? reg_csr_2818 : _GEN_2817; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2819 = 12'hb03 == csr_addr[11:0] ? reg_csr_2819 : _GEN_2818; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2820 = 12'hb04 == csr_addr[11:0] ? reg_csr_2820 : _GEN_2819; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2821 = 12'hb05 == csr_addr[11:0] ? reg_csr_2821 : _GEN_2820; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2822 = 12'hb06 == csr_addr[11:0] ? reg_csr_2822 : _GEN_2821; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2823 = 12'hb07 == csr_addr[11:0] ? reg_csr_2823 : _GEN_2822; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2824 = 12'hb08 == csr_addr[11:0] ? reg_csr_2824 : _GEN_2823; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2825 = 12'hb09 == csr_addr[11:0] ? reg_csr_2825 : _GEN_2824; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2826 = 12'hb0a == csr_addr[11:0] ? reg_csr_2826 : _GEN_2825; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2827 = 12'hb0b == csr_addr[11:0] ? reg_csr_2827 : _GEN_2826; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2828 = 12'hb0c == csr_addr[11:0] ? reg_csr_2828 : _GEN_2827; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2829 = 12'hb0d == csr_addr[11:0] ? reg_csr_2829 : _GEN_2828; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2830 = 12'hb0e == csr_addr[11:0] ? reg_csr_2830 : _GEN_2829; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2831 = 12'hb0f == csr_addr[11:0] ? reg_csr_2831 : _GEN_2830; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2832 = 12'hb10 == csr_addr[11:0] ? reg_csr_2832 : _GEN_2831; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2833 = 12'hb11 == csr_addr[11:0] ? reg_csr_2833 : _GEN_2832; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2834 = 12'hb12 == csr_addr[11:0] ? reg_csr_2834 : _GEN_2833; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2835 = 12'hb13 == csr_addr[11:0] ? reg_csr_2835 : _GEN_2834; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2836 = 12'hb14 == csr_addr[11:0] ? reg_csr_2836 : _GEN_2835; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2837 = 12'hb15 == csr_addr[11:0] ? reg_csr_2837 : _GEN_2836; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2838 = 12'hb16 == csr_addr[11:0] ? reg_csr_2838 : _GEN_2837; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2839 = 12'hb17 == csr_addr[11:0] ? reg_csr_2839 : _GEN_2838; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2840 = 12'hb18 == csr_addr[11:0] ? reg_csr_2840 : _GEN_2839; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2841 = 12'hb19 == csr_addr[11:0] ? reg_csr_2841 : _GEN_2840; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2842 = 12'hb1a == csr_addr[11:0] ? reg_csr_2842 : _GEN_2841; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2843 = 12'hb1b == csr_addr[11:0] ? reg_csr_2843 : _GEN_2842; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2844 = 12'hb1c == csr_addr[11:0] ? reg_csr_2844 : _GEN_2843; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2845 = 12'hb1d == csr_addr[11:0] ? reg_csr_2845 : _GEN_2844; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2846 = 12'hb1e == csr_addr[11:0] ? reg_csr_2846 : _GEN_2845; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2847 = 12'hb1f == csr_addr[11:0] ? reg_csr_2847 : _GEN_2846; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2848 = 12'hb20 == csr_addr[11:0] ? reg_csr_2848 : _GEN_2847; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2849 = 12'hb21 == csr_addr[11:0] ? reg_csr_2849 : _GEN_2848; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2850 = 12'hb22 == csr_addr[11:0] ? reg_csr_2850 : _GEN_2849; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2851 = 12'hb23 == csr_addr[11:0] ? reg_csr_2851 : _GEN_2850; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2852 = 12'hb24 == csr_addr[11:0] ? reg_csr_2852 : _GEN_2851; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2853 = 12'hb25 == csr_addr[11:0] ? reg_csr_2853 : _GEN_2852; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2854 = 12'hb26 == csr_addr[11:0] ? reg_csr_2854 : _GEN_2853; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2855 = 12'hb27 == csr_addr[11:0] ? reg_csr_2855 : _GEN_2854; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2856 = 12'hb28 == csr_addr[11:0] ? reg_csr_2856 : _GEN_2855; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2857 = 12'hb29 == csr_addr[11:0] ? reg_csr_2857 : _GEN_2856; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2858 = 12'hb2a == csr_addr[11:0] ? reg_csr_2858 : _GEN_2857; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2859 = 12'hb2b == csr_addr[11:0] ? reg_csr_2859 : _GEN_2858; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2860 = 12'hb2c == csr_addr[11:0] ? reg_csr_2860 : _GEN_2859; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2861 = 12'hb2d == csr_addr[11:0] ? reg_csr_2861 : _GEN_2860; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2862 = 12'hb2e == csr_addr[11:0] ? reg_csr_2862 : _GEN_2861; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2863 = 12'hb2f == csr_addr[11:0] ? reg_csr_2863 : _GEN_2862; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2864 = 12'hb30 == csr_addr[11:0] ? reg_csr_2864 : _GEN_2863; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2865 = 12'hb31 == csr_addr[11:0] ? reg_csr_2865 : _GEN_2864; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2866 = 12'hb32 == csr_addr[11:0] ? reg_csr_2866 : _GEN_2865; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2867 = 12'hb33 == csr_addr[11:0] ? reg_csr_2867 : _GEN_2866; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2868 = 12'hb34 == csr_addr[11:0] ? reg_csr_2868 : _GEN_2867; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2869 = 12'hb35 == csr_addr[11:0] ? reg_csr_2869 : _GEN_2868; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2870 = 12'hb36 == csr_addr[11:0] ? reg_csr_2870 : _GEN_2869; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2871 = 12'hb37 == csr_addr[11:0] ? reg_csr_2871 : _GEN_2870; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2872 = 12'hb38 == csr_addr[11:0] ? reg_csr_2872 : _GEN_2871; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2873 = 12'hb39 == csr_addr[11:0] ? reg_csr_2873 : _GEN_2872; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2874 = 12'hb3a == csr_addr[11:0] ? reg_csr_2874 : _GEN_2873; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2875 = 12'hb3b == csr_addr[11:0] ? reg_csr_2875 : _GEN_2874; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2876 = 12'hb3c == csr_addr[11:0] ? reg_csr_2876 : _GEN_2875; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2877 = 12'hb3d == csr_addr[11:0] ? reg_csr_2877 : _GEN_2876; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2878 = 12'hb3e == csr_addr[11:0] ? reg_csr_2878 : _GEN_2877; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2879 = 12'hb3f == csr_addr[11:0] ? reg_csr_2879 : _GEN_2878; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2880 = 12'hb40 == csr_addr[11:0] ? reg_csr_2880 : _GEN_2879; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2881 = 12'hb41 == csr_addr[11:0] ? reg_csr_2881 : _GEN_2880; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2882 = 12'hb42 == csr_addr[11:0] ? reg_csr_2882 : _GEN_2881; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2883 = 12'hb43 == csr_addr[11:0] ? reg_csr_2883 : _GEN_2882; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2884 = 12'hb44 == csr_addr[11:0] ? reg_csr_2884 : _GEN_2883; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2885 = 12'hb45 == csr_addr[11:0] ? reg_csr_2885 : _GEN_2884; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2886 = 12'hb46 == csr_addr[11:0] ? reg_csr_2886 : _GEN_2885; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2887 = 12'hb47 == csr_addr[11:0] ? reg_csr_2887 : _GEN_2886; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2888 = 12'hb48 == csr_addr[11:0] ? reg_csr_2888 : _GEN_2887; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2889 = 12'hb49 == csr_addr[11:0] ? reg_csr_2889 : _GEN_2888; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2890 = 12'hb4a == csr_addr[11:0] ? reg_csr_2890 : _GEN_2889; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2891 = 12'hb4b == csr_addr[11:0] ? reg_csr_2891 : _GEN_2890; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2892 = 12'hb4c == csr_addr[11:0] ? reg_csr_2892 : _GEN_2891; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2893 = 12'hb4d == csr_addr[11:0] ? reg_csr_2893 : _GEN_2892; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2894 = 12'hb4e == csr_addr[11:0] ? reg_csr_2894 : _GEN_2893; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2895 = 12'hb4f == csr_addr[11:0] ? reg_csr_2895 : _GEN_2894; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2896 = 12'hb50 == csr_addr[11:0] ? reg_csr_2896 : _GEN_2895; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2897 = 12'hb51 == csr_addr[11:0] ? reg_csr_2897 : _GEN_2896; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2898 = 12'hb52 == csr_addr[11:0] ? reg_csr_2898 : _GEN_2897; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2899 = 12'hb53 == csr_addr[11:0] ? reg_csr_2899 : _GEN_2898; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2900 = 12'hb54 == csr_addr[11:0] ? reg_csr_2900 : _GEN_2899; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2901 = 12'hb55 == csr_addr[11:0] ? reg_csr_2901 : _GEN_2900; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2902 = 12'hb56 == csr_addr[11:0] ? reg_csr_2902 : _GEN_2901; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2903 = 12'hb57 == csr_addr[11:0] ? reg_csr_2903 : _GEN_2902; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2904 = 12'hb58 == csr_addr[11:0] ? reg_csr_2904 : _GEN_2903; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2905 = 12'hb59 == csr_addr[11:0] ? reg_csr_2905 : _GEN_2904; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2906 = 12'hb5a == csr_addr[11:0] ? reg_csr_2906 : _GEN_2905; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2907 = 12'hb5b == csr_addr[11:0] ? reg_csr_2907 : _GEN_2906; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2908 = 12'hb5c == csr_addr[11:0] ? reg_csr_2908 : _GEN_2907; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2909 = 12'hb5d == csr_addr[11:0] ? reg_csr_2909 : _GEN_2908; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2910 = 12'hb5e == csr_addr[11:0] ? reg_csr_2910 : _GEN_2909; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2911 = 12'hb5f == csr_addr[11:0] ? reg_csr_2911 : _GEN_2910; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2912 = 12'hb60 == csr_addr[11:0] ? reg_csr_2912 : _GEN_2911; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2913 = 12'hb61 == csr_addr[11:0] ? reg_csr_2913 : _GEN_2912; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2914 = 12'hb62 == csr_addr[11:0] ? reg_csr_2914 : _GEN_2913; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2915 = 12'hb63 == csr_addr[11:0] ? reg_csr_2915 : _GEN_2914; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2916 = 12'hb64 == csr_addr[11:0] ? reg_csr_2916 : _GEN_2915; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2917 = 12'hb65 == csr_addr[11:0] ? reg_csr_2917 : _GEN_2916; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2918 = 12'hb66 == csr_addr[11:0] ? reg_csr_2918 : _GEN_2917; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2919 = 12'hb67 == csr_addr[11:0] ? reg_csr_2919 : _GEN_2918; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2920 = 12'hb68 == csr_addr[11:0] ? reg_csr_2920 : _GEN_2919; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2921 = 12'hb69 == csr_addr[11:0] ? reg_csr_2921 : _GEN_2920; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2922 = 12'hb6a == csr_addr[11:0] ? reg_csr_2922 : _GEN_2921; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2923 = 12'hb6b == csr_addr[11:0] ? reg_csr_2923 : _GEN_2922; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2924 = 12'hb6c == csr_addr[11:0] ? reg_csr_2924 : _GEN_2923; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2925 = 12'hb6d == csr_addr[11:0] ? reg_csr_2925 : _GEN_2924; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2926 = 12'hb6e == csr_addr[11:0] ? reg_csr_2926 : _GEN_2925; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2927 = 12'hb6f == csr_addr[11:0] ? reg_csr_2927 : _GEN_2926; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2928 = 12'hb70 == csr_addr[11:0] ? reg_csr_2928 : _GEN_2927; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2929 = 12'hb71 == csr_addr[11:0] ? reg_csr_2929 : _GEN_2928; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2930 = 12'hb72 == csr_addr[11:0] ? reg_csr_2930 : _GEN_2929; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2931 = 12'hb73 == csr_addr[11:0] ? reg_csr_2931 : _GEN_2930; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2932 = 12'hb74 == csr_addr[11:0] ? reg_csr_2932 : _GEN_2931; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2933 = 12'hb75 == csr_addr[11:0] ? reg_csr_2933 : _GEN_2932; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2934 = 12'hb76 == csr_addr[11:0] ? reg_csr_2934 : _GEN_2933; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2935 = 12'hb77 == csr_addr[11:0] ? reg_csr_2935 : _GEN_2934; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2936 = 12'hb78 == csr_addr[11:0] ? reg_csr_2936 : _GEN_2935; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2937 = 12'hb79 == csr_addr[11:0] ? reg_csr_2937 : _GEN_2936; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2938 = 12'hb7a == csr_addr[11:0] ? reg_csr_2938 : _GEN_2937; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2939 = 12'hb7b == csr_addr[11:0] ? reg_csr_2939 : _GEN_2938; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2940 = 12'hb7c == csr_addr[11:0] ? reg_csr_2940 : _GEN_2939; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2941 = 12'hb7d == csr_addr[11:0] ? reg_csr_2941 : _GEN_2940; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2942 = 12'hb7e == csr_addr[11:0] ? reg_csr_2942 : _GEN_2941; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2943 = 12'hb7f == csr_addr[11:0] ? reg_csr_2943 : _GEN_2942; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2944 = 12'hb80 == csr_addr[11:0] ? reg_csr_2944 : _GEN_2943; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2945 = 12'hb81 == csr_addr[11:0] ? reg_csr_2945 : _GEN_2944; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2946 = 12'hb82 == csr_addr[11:0] ? reg_csr_2946 : _GEN_2945; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2947 = 12'hb83 == csr_addr[11:0] ? reg_csr_2947 : _GEN_2946; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2948 = 12'hb84 == csr_addr[11:0] ? reg_csr_2948 : _GEN_2947; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2949 = 12'hb85 == csr_addr[11:0] ? reg_csr_2949 : _GEN_2948; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2950 = 12'hb86 == csr_addr[11:0] ? reg_csr_2950 : _GEN_2949; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2951 = 12'hb87 == csr_addr[11:0] ? reg_csr_2951 : _GEN_2950; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2952 = 12'hb88 == csr_addr[11:0] ? reg_csr_2952 : _GEN_2951; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2953 = 12'hb89 == csr_addr[11:0] ? reg_csr_2953 : _GEN_2952; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2954 = 12'hb8a == csr_addr[11:0] ? reg_csr_2954 : _GEN_2953; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2955 = 12'hb8b == csr_addr[11:0] ? reg_csr_2955 : _GEN_2954; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2956 = 12'hb8c == csr_addr[11:0] ? reg_csr_2956 : _GEN_2955; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2957 = 12'hb8d == csr_addr[11:0] ? reg_csr_2957 : _GEN_2956; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2958 = 12'hb8e == csr_addr[11:0] ? reg_csr_2958 : _GEN_2957; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2959 = 12'hb8f == csr_addr[11:0] ? reg_csr_2959 : _GEN_2958; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2960 = 12'hb90 == csr_addr[11:0] ? reg_csr_2960 : _GEN_2959; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2961 = 12'hb91 == csr_addr[11:0] ? reg_csr_2961 : _GEN_2960; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2962 = 12'hb92 == csr_addr[11:0] ? reg_csr_2962 : _GEN_2961; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2963 = 12'hb93 == csr_addr[11:0] ? reg_csr_2963 : _GEN_2962; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2964 = 12'hb94 == csr_addr[11:0] ? reg_csr_2964 : _GEN_2963; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2965 = 12'hb95 == csr_addr[11:0] ? reg_csr_2965 : _GEN_2964; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2966 = 12'hb96 == csr_addr[11:0] ? reg_csr_2966 : _GEN_2965; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2967 = 12'hb97 == csr_addr[11:0] ? reg_csr_2967 : _GEN_2966; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2968 = 12'hb98 == csr_addr[11:0] ? reg_csr_2968 : _GEN_2967; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2969 = 12'hb99 == csr_addr[11:0] ? reg_csr_2969 : _GEN_2968; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2970 = 12'hb9a == csr_addr[11:0] ? reg_csr_2970 : _GEN_2969; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2971 = 12'hb9b == csr_addr[11:0] ? reg_csr_2971 : _GEN_2970; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2972 = 12'hb9c == csr_addr[11:0] ? reg_csr_2972 : _GEN_2971; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2973 = 12'hb9d == csr_addr[11:0] ? reg_csr_2973 : _GEN_2972; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2974 = 12'hb9e == csr_addr[11:0] ? reg_csr_2974 : _GEN_2973; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2975 = 12'hb9f == csr_addr[11:0] ? reg_csr_2975 : _GEN_2974; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2976 = 12'hba0 == csr_addr[11:0] ? reg_csr_2976 : _GEN_2975; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2977 = 12'hba1 == csr_addr[11:0] ? reg_csr_2977 : _GEN_2976; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2978 = 12'hba2 == csr_addr[11:0] ? reg_csr_2978 : _GEN_2977; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2979 = 12'hba3 == csr_addr[11:0] ? reg_csr_2979 : _GEN_2978; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2980 = 12'hba4 == csr_addr[11:0] ? reg_csr_2980 : _GEN_2979; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2981 = 12'hba5 == csr_addr[11:0] ? reg_csr_2981 : _GEN_2980; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2982 = 12'hba6 == csr_addr[11:0] ? reg_csr_2982 : _GEN_2981; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2983 = 12'hba7 == csr_addr[11:0] ? reg_csr_2983 : _GEN_2982; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2984 = 12'hba8 == csr_addr[11:0] ? reg_csr_2984 : _GEN_2983; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2985 = 12'hba9 == csr_addr[11:0] ? reg_csr_2985 : _GEN_2984; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2986 = 12'hbaa == csr_addr[11:0] ? reg_csr_2986 : _GEN_2985; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2987 = 12'hbab == csr_addr[11:0] ? reg_csr_2987 : _GEN_2986; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2988 = 12'hbac == csr_addr[11:0] ? reg_csr_2988 : _GEN_2987; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2989 = 12'hbad == csr_addr[11:0] ? reg_csr_2989 : _GEN_2988; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2990 = 12'hbae == csr_addr[11:0] ? reg_csr_2990 : _GEN_2989; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2991 = 12'hbaf == csr_addr[11:0] ? reg_csr_2991 : _GEN_2990; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2992 = 12'hbb0 == csr_addr[11:0] ? reg_csr_2992 : _GEN_2991; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2993 = 12'hbb1 == csr_addr[11:0] ? reg_csr_2993 : _GEN_2992; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2994 = 12'hbb2 == csr_addr[11:0] ? reg_csr_2994 : _GEN_2993; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2995 = 12'hbb3 == csr_addr[11:0] ? reg_csr_2995 : _GEN_2994; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2996 = 12'hbb4 == csr_addr[11:0] ? reg_csr_2996 : _GEN_2995; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2997 = 12'hbb5 == csr_addr[11:0] ? reg_csr_2997 : _GEN_2996; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2998 = 12'hbb6 == csr_addr[11:0] ? reg_csr_2998 : _GEN_2997; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_2999 = 12'hbb7 == csr_addr[11:0] ? reg_csr_2999 : _GEN_2998; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3000 = 12'hbb8 == csr_addr[11:0] ? reg_csr_3000 : _GEN_2999; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3001 = 12'hbb9 == csr_addr[11:0] ? reg_csr_3001 : _GEN_3000; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3002 = 12'hbba == csr_addr[11:0] ? reg_csr_3002 : _GEN_3001; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3003 = 12'hbbb == csr_addr[11:0] ? reg_csr_3003 : _GEN_3002; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3004 = 12'hbbc == csr_addr[11:0] ? reg_csr_3004 : _GEN_3003; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3005 = 12'hbbd == csr_addr[11:0] ? reg_csr_3005 : _GEN_3004; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3006 = 12'hbbe == csr_addr[11:0] ? reg_csr_3006 : _GEN_3005; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3007 = 12'hbbf == csr_addr[11:0] ? reg_csr_3007 : _GEN_3006; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3008 = 12'hbc0 == csr_addr[11:0] ? reg_csr_3008 : _GEN_3007; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3009 = 12'hbc1 == csr_addr[11:0] ? reg_csr_3009 : _GEN_3008; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3010 = 12'hbc2 == csr_addr[11:0] ? reg_csr_3010 : _GEN_3009; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3011 = 12'hbc3 == csr_addr[11:0] ? reg_csr_3011 : _GEN_3010; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3012 = 12'hbc4 == csr_addr[11:0] ? reg_csr_3012 : _GEN_3011; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3013 = 12'hbc5 == csr_addr[11:0] ? reg_csr_3013 : _GEN_3012; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3014 = 12'hbc6 == csr_addr[11:0] ? reg_csr_3014 : _GEN_3013; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3015 = 12'hbc7 == csr_addr[11:0] ? reg_csr_3015 : _GEN_3014; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3016 = 12'hbc8 == csr_addr[11:0] ? reg_csr_3016 : _GEN_3015; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3017 = 12'hbc9 == csr_addr[11:0] ? reg_csr_3017 : _GEN_3016; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3018 = 12'hbca == csr_addr[11:0] ? reg_csr_3018 : _GEN_3017; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3019 = 12'hbcb == csr_addr[11:0] ? reg_csr_3019 : _GEN_3018; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3020 = 12'hbcc == csr_addr[11:0] ? reg_csr_3020 : _GEN_3019; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3021 = 12'hbcd == csr_addr[11:0] ? reg_csr_3021 : _GEN_3020; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3022 = 12'hbce == csr_addr[11:0] ? reg_csr_3022 : _GEN_3021; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3023 = 12'hbcf == csr_addr[11:0] ? reg_csr_3023 : _GEN_3022; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3024 = 12'hbd0 == csr_addr[11:0] ? reg_csr_3024 : _GEN_3023; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3025 = 12'hbd1 == csr_addr[11:0] ? reg_csr_3025 : _GEN_3024; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3026 = 12'hbd2 == csr_addr[11:0] ? reg_csr_3026 : _GEN_3025; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3027 = 12'hbd3 == csr_addr[11:0] ? reg_csr_3027 : _GEN_3026; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3028 = 12'hbd4 == csr_addr[11:0] ? reg_csr_3028 : _GEN_3027; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3029 = 12'hbd5 == csr_addr[11:0] ? reg_csr_3029 : _GEN_3028; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3030 = 12'hbd6 == csr_addr[11:0] ? reg_csr_3030 : _GEN_3029; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3031 = 12'hbd7 == csr_addr[11:0] ? reg_csr_3031 : _GEN_3030; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3032 = 12'hbd8 == csr_addr[11:0] ? reg_csr_3032 : _GEN_3031; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3033 = 12'hbd9 == csr_addr[11:0] ? reg_csr_3033 : _GEN_3032; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3034 = 12'hbda == csr_addr[11:0] ? reg_csr_3034 : _GEN_3033; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3035 = 12'hbdb == csr_addr[11:0] ? reg_csr_3035 : _GEN_3034; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3036 = 12'hbdc == csr_addr[11:0] ? reg_csr_3036 : _GEN_3035; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3037 = 12'hbdd == csr_addr[11:0] ? reg_csr_3037 : _GEN_3036; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3038 = 12'hbde == csr_addr[11:0] ? reg_csr_3038 : _GEN_3037; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3039 = 12'hbdf == csr_addr[11:0] ? reg_csr_3039 : _GEN_3038; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3040 = 12'hbe0 == csr_addr[11:0] ? reg_csr_3040 : _GEN_3039; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3041 = 12'hbe1 == csr_addr[11:0] ? reg_csr_3041 : _GEN_3040; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3042 = 12'hbe2 == csr_addr[11:0] ? reg_csr_3042 : _GEN_3041; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3043 = 12'hbe3 == csr_addr[11:0] ? reg_csr_3043 : _GEN_3042; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3044 = 12'hbe4 == csr_addr[11:0] ? reg_csr_3044 : _GEN_3043; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3045 = 12'hbe5 == csr_addr[11:0] ? reg_csr_3045 : _GEN_3044; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3046 = 12'hbe6 == csr_addr[11:0] ? reg_csr_3046 : _GEN_3045; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3047 = 12'hbe7 == csr_addr[11:0] ? reg_csr_3047 : _GEN_3046; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3048 = 12'hbe8 == csr_addr[11:0] ? reg_csr_3048 : _GEN_3047; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3049 = 12'hbe9 == csr_addr[11:0] ? reg_csr_3049 : _GEN_3048; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3050 = 12'hbea == csr_addr[11:0] ? reg_csr_3050 : _GEN_3049; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3051 = 12'hbeb == csr_addr[11:0] ? reg_csr_3051 : _GEN_3050; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3052 = 12'hbec == csr_addr[11:0] ? reg_csr_3052 : _GEN_3051; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3053 = 12'hbed == csr_addr[11:0] ? reg_csr_3053 : _GEN_3052; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3054 = 12'hbee == csr_addr[11:0] ? reg_csr_3054 : _GEN_3053; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3055 = 12'hbef == csr_addr[11:0] ? reg_csr_3055 : _GEN_3054; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3056 = 12'hbf0 == csr_addr[11:0] ? reg_csr_3056 : _GEN_3055; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3057 = 12'hbf1 == csr_addr[11:0] ? reg_csr_3057 : _GEN_3056; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3058 = 12'hbf2 == csr_addr[11:0] ? reg_csr_3058 : _GEN_3057; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3059 = 12'hbf3 == csr_addr[11:0] ? reg_csr_3059 : _GEN_3058; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3060 = 12'hbf4 == csr_addr[11:0] ? reg_csr_3060 : _GEN_3059; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3061 = 12'hbf5 == csr_addr[11:0] ? reg_csr_3061 : _GEN_3060; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3062 = 12'hbf6 == csr_addr[11:0] ? reg_csr_3062 : _GEN_3061; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3063 = 12'hbf7 == csr_addr[11:0] ? reg_csr_3063 : _GEN_3062; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3064 = 12'hbf8 == csr_addr[11:0] ? reg_csr_3064 : _GEN_3063; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3065 = 12'hbf9 == csr_addr[11:0] ? reg_csr_3065 : _GEN_3064; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3066 = 12'hbfa == csr_addr[11:0] ? reg_csr_3066 : _GEN_3065; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3067 = 12'hbfb == csr_addr[11:0] ? reg_csr_3067 : _GEN_3066; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3068 = 12'hbfc == csr_addr[11:0] ? reg_csr_3068 : _GEN_3067; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3069 = 12'hbfd == csr_addr[11:0] ? reg_csr_3069 : _GEN_3068; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3070 = 12'hbfe == csr_addr[11:0] ? reg_csr_3070 : _GEN_3069; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3071 = 12'hbff == csr_addr[11:0] ? reg_csr_3071 : _GEN_3070; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3072 = 12'hc00 == csr_addr[11:0] ? reg_csr_3072 : _GEN_3071; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3073 = 12'hc01 == csr_addr[11:0] ? reg_csr_3073 : _GEN_3072; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3074 = 12'hc02 == csr_addr[11:0] ? reg_csr_3074 : _GEN_3073; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3075 = 12'hc03 == csr_addr[11:0] ? reg_csr_3075 : _GEN_3074; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3076 = 12'hc04 == csr_addr[11:0] ? reg_csr_3076 : _GEN_3075; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3077 = 12'hc05 == csr_addr[11:0] ? reg_csr_3077 : _GEN_3076; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3078 = 12'hc06 == csr_addr[11:0] ? reg_csr_3078 : _GEN_3077; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3079 = 12'hc07 == csr_addr[11:0] ? reg_csr_3079 : _GEN_3078; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3080 = 12'hc08 == csr_addr[11:0] ? reg_csr_3080 : _GEN_3079; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3081 = 12'hc09 == csr_addr[11:0] ? reg_csr_3081 : _GEN_3080; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3082 = 12'hc0a == csr_addr[11:0] ? reg_csr_3082 : _GEN_3081; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3083 = 12'hc0b == csr_addr[11:0] ? reg_csr_3083 : _GEN_3082; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3084 = 12'hc0c == csr_addr[11:0] ? reg_csr_3084 : _GEN_3083; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3085 = 12'hc0d == csr_addr[11:0] ? reg_csr_3085 : _GEN_3084; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3086 = 12'hc0e == csr_addr[11:0] ? reg_csr_3086 : _GEN_3085; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3087 = 12'hc0f == csr_addr[11:0] ? reg_csr_3087 : _GEN_3086; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3088 = 12'hc10 == csr_addr[11:0] ? reg_csr_3088 : _GEN_3087; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3089 = 12'hc11 == csr_addr[11:0] ? reg_csr_3089 : _GEN_3088; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3090 = 12'hc12 == csr_addr[11:0] ? reg_csr_3090 : _GEN_3089; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3091 = 12'hc13 == csr_addr[11:0] ? reg_csr_3091 : _GEN_3090; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3092 = 12'hc14 == csr_addr[11:0] ? reg_csr_3092 : _GEN_3091; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3093 = 12'hc15 == csr_addr[11:0] ? reg_csr_3093 : _GEN_3092; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3094 = 12'hc16 == csr_addr[11:0] ? reg_csr_3094 : _GEN_3093; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3095 = 12'hc17 == csr_addr[11:0] ? reg_csr_3095 : _GEN_3094; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3096 = 12'hc18 == csr_addr[11:0] ? reg_csr_3096 : _GEN_3095; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3097 = 12'hc19 == csr_addr[11:0] ? reg_csr_3097 : _GEN_3096; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3098 = 12'hc1a == csr_addr[11:0] ? reg_csr_3098 : _GEN_3097; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3099 = 12'hc1b == csr_addr[11:0] ? reg_csr_3099 : _GEN_3098; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3100 = 12'hc1c == csr_addr[11:0] ? reg_csr_3100 : _GEN_3099; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3101 = 12'hc1d == csr_addr[11:0] ? reg_csr_3101 : _GEN_3100; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3102 = 12'hc1e == csr_addr[11:0] ? reg_csr_3102 : _GEN_3101; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3103 = 12'hc1f == csr_addr[11:0] ? reg_csr_3103 : _GEN_3102; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3104 = 12'hc20 == csr_addr[11:0] ? reg_csr_3104 : _GEN_3103; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3105 = 12'hc21 == csr_addr[11:0] ? reg_csr_3105 : _GEN_3104; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3106 = 12'hc22 == csr_addr[11:0] ? reg_csr_3106 : _GEN_3105; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3107 = 12'hc23 == csr_addr[11:0] ? reg_csr_3107 : _GEN_3106; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3108 = 12'hc24 == csr_addr[11:0] ? reg_csr_3108 : _GEN_3107; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3109 = 12'hc25 == csr_addr[11:0] ? reg_csr_3109 : _GEN_3108; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3110 = 12'hc26 == csr_addr[11:0] ? reg_csr_3110 : _GEN_3109; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3111 = 12'hc27 == csr_addr[11:0] ? reg_csr_3111 : _GEN_3110; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3112 = 12'hc28 == csr_addr[11:0] ? reg_csr_3112 : _GEN_3111; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3113 = 12'hc29 == csr_addr[11:0] ? reg_csr_3113 : _GEN_3112; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3114 = 12'hc2a == csr_addr[11:0] ? reg_csr_3114 : _GEN_3113; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3115 = 12'hc2b == csr_addr[11:0] ? reg_csr_3115 : _GEN_3114; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3116 = 12'hc2c == csr_addr[11:0] ? reg_csr_3116 : _GEN_3115; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3117 = 12'hc2d == csr_addr[11:0] ? reg_csr_3117 : _GEN_3116; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3118 = 12'hc2e == csr_addr[11:0] ? reg_csr_3118 : _GEN_3117; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3119 = 12'hc2f == csr_addr[11:0] ? reg_csr_3119 : _GEN_3118; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3120 = 12'hc30 == csr_addr[11:0] ? reg_csr_3120 : _GEN_3119; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3121 = 12'hc31 == csr_addr[11:0] ? reg_csr_3121 : _GEN_3120; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3122 = 12'hc32 == csr_addr[11:0] ? reg_csr_3122 : _GEN_3121; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3123 = 12'hc33 == csr_addr[11:0] ? reg_csr_3123 : _GEN_3122; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3124 = 12'hc34 == csr_addr[11:0] ? reg_csr_3124 : _GEN_3123; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3125 = 12'hc35 == csr_addr[11:0] ? reg_csr_3125 : _GEN_3124; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3126 = 12'hc36 == csr_addr[11:0] ? reg_csr_3126 : _GEN_3125; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3127 = 12'hc37 == csr_addr[11:0] ? reg_csr_3127 : _GEN_3126; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3128 = 12'hc38 == csr_addr[11:0] ? reg_csr_3128 : _GEN_3127; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3129 = 12'hc39 == csr_addr[11:0] ? reg_csr_3129 : _GEN_3128; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3130 = 12'hc3a == csr_addr[11:0] ? reg_csr_3130 : _GEN_3129; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3131 = 12'hc3b == csr_addr[11:0] ? reg_csr_3131 : _GEN_3130; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3132 = 12'hc3c == csr_addr[11:0] ? reg_csr_3132 : _GEN_3131; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3133 = 12'hc3d == csr_addr[11:0] ? reg_csr_3133 : _GEN_3132; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3134 = 12'hc3e == csr_addr[11:0] ? reg_csr_3134 : _GEN_3133; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3135 = 12'hc3f == csr_addr[11:0] ? reg_csr_3135 : _GEN_3134; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3136 = 12'hc40 == csr_addr[11:0] ? reg_csr_3136 : _GEN_3135; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3137 = 12'hc41 == csr_addr[11:0] ? reg_csr_3137 : _GEN_3136; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3138 = 12'hc42 == csr_addr[11:0] ? reg_csr_3138 : _GEN_3137; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3139 = 12'hc43 == csr_addr[11:0] ? reg_csr_3139 : _GEN_3138; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3140 = 12'hc44 == csr_addr[11:0] ? reg_csr_3140 : _GEN_3139; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3141 = 12'hc45 == csr_addr[11:0] ? reg_csr_3141 : _GEN_3140; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3142 = 12'hc46 == csr_addr[11:0] ? reg_csr_3142 : _GEN_3141; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3143 = 12'hc47 == csr_addr[11:0] ? reg_csr_3143 : _GEN_3142; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3144 = 12'hc48 == csr_addr[11:0] ? reg_csr_3144 : _GEN_3143; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3145 = 12'hc49 == csr_addr[11:0] ? reg_csr_3145 : _GEN_3144; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3146 = 12'hc4a == csr_addr[11:0] ? reg_csr_3146 : _GEN_3145; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3147 = 12'hc4b == csr_addr[11:0] ? reg_csr_3147 : _GEN_3146; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3148 = 12'hc4c == csr_addr[11:0] ? reg_csr_3148 : _GEN_3147; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3149 = 12'hc4d == csr_addr[11:0] ? reg_csr_3149 : _GEN_3148; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3150 = 12'hc4e == csr_addr[11:0] ? reg_csr_3150 : _GEN_3149; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3151 = 12'hc4f == csr_addr[11:0] ? reg_csr_3151 : _GEN_3150; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3152 = 12'hc50 == csr_addr[11:0] ? reg_csr_3152 : _GEN_3151; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3153 = 12'hc51 == csr_addr[11:0] ? reg_csr_3153 : _GEN_3152; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3154 = 12'hc52 == csr_addr[11:0] ? reg_csr_3154 : _GEN_3153; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3155 = 12'hc53 == csr_addr[11:0] ? reg_csr_3155 : _GEN_3154; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3156 = 12'hc54 == csr_addr[11:0] ? reg_csr_3156 : _GEN_3155; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3157 = 12'hc55 == csr_addr[11:0] ? reg_csr_3157 : _GEN_3156; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3158 = 12'hc56 == csr_addr[11:0] ? reg_csr_3158 : _GEN_3157; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3159 = 12'hc57 == csr_addr[11:0] ? reg_csr_3159 : _GEN_3158; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3160 = 12'hc58 == csr_addr[11:0] ? reg_csr_3160 : _GEN_3159; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3161 = 12'hc59 == csr_addr[11:0] ? reg_csr_3161 : _GEN_3160; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3162 = 12'hc5a == csr_addr[11:0] ? reg_csr_3162 : _GEN_3161; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3163 = 12'hc5b == csr_addr[11:0] ? reg_csr_3163 : _GEN_3162; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3164 = 12'hc5c == csr_addr[11:0] ? reg_csr_3164 : _GEN_3163; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3165 = 12'hc5d == csr_addr[11:0] ? reg_csr_3165 : _GEN_3164; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3166 = 12'hc5e == csr_addr[11:0] ? reg_csr_3166 : _GEN_3165; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3167 = 12'hc5f == csr_addr[11:0] ? reg_csr_3167 : _GEN_3166; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3168 = 12'hc60 == csr_addr[11:0] ? reg_csr_3168 : _GEN_3167; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3169 = 12'hc61 == csr_addr[11:0] ? reg_csr_3169 : _GEN_3168; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3170 = 12'hc62 == csr_addr[11:0] ? reg_csr_3170 : _GEN_3169; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3171 = 12'hc63 == csr_addr[11:0] ? reg_csr_3171 : _GEN_3170; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3172 = 12'hc64 == csr_addr[11:0] ? reg_csr_3172 : _GEN_3171; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3173 = 12'hc65 == csr_addr[11:0] ? reg_csr_3173 : _GEN_3172; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3174 = 12'hc66 == csr_addr[11:0] ? reg_csr_3174 : _GEN_3173; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3175 = 12'hc67 == csr_addr[11:0] ? reg_csr_3175 : _GEN_3174; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3176 = 12'hc68 == csr_addr[11:0] ? reg_csr_3176 : _GEN_3175; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3177 = 12'hc69 == csr_addr[11:0] ? reg_csr_3177 : _GEN_3176; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3178 = 12'hc6a == csr_addr[11:0] ? reg_csr_3178 : _GEN_3177; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3179 = 12'hc6b == csr_addr[11:0] ? reg_csr_3179 : _GEN_3178; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3180 = 12'hc6c == csr_addr[11:0] ? reg_csr_3180 : _GEN_3179; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3181 = 12'hc6d == csr_addr[11:0] ? reg_csr_3181 : _GEN_3180; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3182 = 12'hc6e == csr_addr[11:0] ? reg_csr_3182 : _GEN_3181; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3183 = 12'hc6f == csr_addr[11:0] ? reg_csr_3183 : _GEN_3182; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3184 = 12'hc70 == csr_addr[11:0] ? reg_csr_3184 : _GEN_3183; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3185 = 12'hc71 == csr_addr[11:0] ? reg_csr_3185 : _GEN_3184; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3186 = 12'hc72 == csr_addr[11:0] ? reg_csr_3186 : _GEN_3185; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3187 = 12'hc73 == csr_addr[11:0] ? reg_csr_3187 : _GEN_3186; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3188 = 12'hc74 == csr_addr[11:0] ? reg_csr_3188 : _GEN_3187; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3189 = 12'hc75 == csr_addr[11:0] ? reg_csr_3189 : _GEN_3188; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3190 = 12'hc76 == csr_addr[11:0] ? reg_csr_3190 : _GEN_3189; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3191 = 12'hc77 == csr_addr[11:0] ? reg_csr_3191 : _GEN_3190; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3192 = 12'hc78 == csr_addr[11:0] ? reg_csr_3192 : _GEN_3191; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3193 = 12'hc79 == csr_addr[11:0] ? reg_csr_3193 : _GEN_3192; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3194 = 12'hc7a == csr_addr[11:0] ? reg_csr_3194 : _GEN_3193; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3195 = 12'hc7b == csr_addr[11:0] ? reg_csr_3195 : _GEN_3194; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3196 = 12'hc7c == csr_addr[11:0] ? reg_csr_3196 : _GEN_3195; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3197 = 12'hc7d == csr_addr[11:0] ? reg_csr_3197 : _GEN_3196; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3198 = 12'hc7e == csr_addr[11:0] ? reg_csr_3198 : _GEN_3197; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3199 = 12'hc7f == csr_addr[11:0] ? reg_csr_3199 : _GEN_3198; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3200 = 12'hc80 == csr_addr[11:0] ? reg_csr_3200 : _GEN_3199; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3201 = 12'hc81 == csr_addr[11:0] ? reg_csr_3201 : _GEN_3200; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3202 = 12'hc82 == csr_addr[11:0] ? reg_csr_3202 : _GEN_3201; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3203 = 12'hc83 == csr_addr[11:0] ? reg_csr_3203 : _GEN_3202; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3204 = 12'hc84 == csr_addr[11:0] ? reg_csr_3204 : _GEN_3203; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3205 = 12'hc85 == csr_addr[11:0] ? reg_csr_3205 : _GEN_3204; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3206 = 12'hc86 == csr_addr[11:0] ? reg_csr_3206 : _GEN_3205; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3207 = 12'hc87 == csr_addr[11:0] ? reg_csr_3207 : _GEN_3206; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3208 = 12'hc88 == csr_addr[11:0] ? reg_csr_3208 : _GEN_3207; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3209 = 12'hc89 == csr_addr[11:0] ? reg_csr_3209 : _GEN_3208; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3210 = 12'hc8a == csr_addr[11:0] ? reg_csr_3210 : _GEN_3209; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3211 = 12'hc8b == csr_addr[11:0] ? reg_csr_3211 : _GEN_3210; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3212 = 12'hc8c == csr_addr[11:0] ? reg_csr_3212 : _GEN_3211; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3213 = 12'hc8d == csr_addr[11:0] ? reg_csr_3213 : _GEN_3212; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3214 = 12'hc8e == csr_addr[11:0] ? reg_csr_3214 : _GEN_3213; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3215 = 12'hc8f == csr_addr[11:0] ? reg_csr_3215 : _GEN_3214; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3216 = 12'hc90 == csr_addr[11:0] ? reg_csr_3216 : _GEN_3215; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3217 = 12'hc91 == csr_addr[11:0] ? reg_csr_3217 : _GEN_3216; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3218 = 12'hc92 == csr_addr[11:0] ? reg_csr_3218 : _GEN_3217; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3219 = 12'hc93 == csr_addr[11:0] ? reg_csr_3219 : _GEN_3218; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3220 = 12'hc94 == csr_addr[11:0] ? reg_csr_3220 : _GEN_3219; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3221 = 12'hc95 == csr_addr[11:0] ? reg_csr_3221 : _GEN_3220; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3222 = 12'hc96 == csr_addr[11:0] ? reg_csr_3222 : _GEN_3221; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3223 = 12'hc97 == csr_addr[11:0] ? reg_csr_3223 : _GEN_3222; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3224 = 12'hc98 == csr_addr[11:0] ? reg_csr_3224 : _GEN_3223; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3225 = 12'hc99 == csr_addr[11:0] ? reg_csr_3225 : _GEN_3224; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3226 = 12'hc9a == csr_addr[11:0] ? reg_csr_3226 : _GEN_3225; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3227 = 12'hc9b == csr_addr[11:0] ? reg_csr_3227 : _GEN_3226; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3228 = 12'hc9c == csr_addr[11:0] ? reg_csr_3228 : _GEN_3227; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3229 = 12'hc9d == csr_addr[11:0] ? reg_csr_3229 : _GEN_3228; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3230 = 12'hc9e == csr_addr[11:0] ? reg_csr_3230 : _GEN_3229; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3231 = 12'hc9f == csr_addr[11:0] ? reg_csr_3231 : _GEN_3230; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3232 = 12'hca0 == csr_addr[11:0] ? reg_csr_3232 : _GEN_3231; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3233 = 12'hca1 == csr_addr[11:0] ? reg_csr_3233 : _GEN_3232; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3234 = 12'hca2 == csr_addr[11:0] ? reg_csr_3234 : _GEN_3233; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3235 = 12'hca3 == csr_addr[11:0] ? reg_csr_3235 : _GEN_3234; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3236 = 12'hca4 == csr_addr[11:0] ? reg_csr_3236 : _GEN_3235; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3237 = 12'hca5 == csr_addr[11:0] ? reg_csr_3237 : _GEN_3236; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3238 = 12'hca6 == csr_addr[11:0] ? reg_csr_3238 : _GEN_3237; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3239 = 12'hca7 == csr_addr[11:0] ? reg_csr_3239 : _GEN_3238; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3240 = 12'hca8 == csr_addr[11:0] ? reg_csr_3240 : _GEN_3239; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3241 = 12'hca9 == csr_addr[11:0] ? reg_csr_3241 : _GEN_3240; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3242 = 12'hcaa == csr_addr[11:0] ? reg_csr_3242 : _GEN_3241; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3243 = 12'hcab == csr_addr[11:0] ? reg_csr_3243 : _GEN_3242; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3244 = 12'hcac == csr_addr[11:0] ? reg_csr_3244 : _GEN_3243; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3245 = 12'hcad == csr_addr[11:0] ? reg_csr_3245 : _GEN_3244; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3246 = 12'hcae == csr_addr[11:0] ? reg_csr_3246 : _GEN_3245; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3247 = 12'hcaf == csr_addr[11:0] ? reg_csr_3247 : _GEN_3246; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3248 = 12'hcb0 == csr_addr[11:0] ? reg_csr_3248 : _GEN_3247; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3249 = 12'hcb1 == csr_addr[11:0] ? reg_csr_3249 : _GEN_3248; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3250 = 12'hcb2 == csr_addr[11:0] ? reg_csr_3250 : _GEN_3249; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3251 = 12'hcb3 == csr_addr[11:0] ? reg_csr_3251 : _GEN_3250; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3252 = 12'hcb4 == csr_addr[11:0] ? reg_csr_3252 : _GEN_3251; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3253 = 12'hcb5 == csr_addr[11:0] ? reg_csr_3253 : _GEN_3252; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3254 = 12'hcb6 == csr_addr[11:0] ? reg_csr_3254 : _GEN_3253; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3255 = 12'hcb7 == csr_addr[11:0] ? reg_csr_3255 : _GEN_3254; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3256 = 12'hcb8 == csr_addr[11:0] ? reg_csr_3256 : _GEN_3255; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3257 = 12'hcb9 == csr_addr[11:0] ? reg_csr_3257 : _GEN_3256; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3258 = 12'hcba == csr_addr[11:0] ? reg_csr_3258 : _GEN_3257; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3259 = 12'hcbb == csr_addr[11:0] ? reg_csr_3259 : _GEN_3258; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3260 = 12'hcbc == csr_addr[11:0] ? reg_csr_3260 : _GEN_3259; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3261 = 12'hcbd == csr_addr[11:0] ? reg_csr_3261 : _GEN_3260; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3262 = 12'hcbe == csr_addr[11:0] ? reg_csr_3262 : _GEN_3261; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3263 = 12'hcbf == csr_addr[11:0] ? reg_csr_3263 : _GEN_3262; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3264 = 12'hcc0 == csr_addr[11:0] ? reg_csr_3264 : _GEN_3263; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3265 = 12'hcc1 == csr_addr[11:0] ? reg_csr_3265 : _GEN_3264; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3266 = 12'hcc2 == csr_addr[11:0] ? reg_csr_3266 : _GEN_3265; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3267 = 12'hcc3 == csr_addr[11:0] ? reg_csr_3267 : _GEN_3266; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3268 = 12'hcc4 == csr_addr[11:0] ? reg_csr_3268 : _GEN_3267; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3269 = 12'hcc5 == csr_addr[11:0] ? reg_csr_3269 : _GEN_3268; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3270 = 12'hcc6 == csr_addr[11:0] ? reg_csr_3270 : _GEN_3269; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3271 = 12'hcc7 == csr_addr[11:0] ? reg_csr_3271 : _GEN_3270; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3272 = 12'hcc8 == csr_addr[11:0] ? reg_csr_3272 : _GEN_3271; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3273 = 12'hcc9 == csr_addr[11:0] ? reg_csr_3273 : _GEN_3272; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3274 = 12'hcca == csr_addr[11:0] ? reg_csr_3274 : _GEN_3273; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3275 = 12'hccb == csr_addr[11:0] ? reg_csr_3275 : _GEN_3274; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3276 = 12'hccc == csr_addr[11:0] ? reg_csr_3276 : _GEN_3275; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3277 = 12'hccd == csr_addr[11:0] ? reg_csr_3277 : _GEN_3276; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3278 = 12'hcce == csr_addr[11:0] ? reg_csr_3278 : _GEN_3277; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3279 = 12'hccf == csr_addr[11:0] ? reg_csr_3279 : _GEN_3278; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3280 = 12'hcd0 == csr_addr[11:0] ? reg_csr_3280 : _GEN_3279; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3281 = 12'hcd1 == csr_addr[11:0] ? reg_csr_3281 : _GEN_3280; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3282 = 12'hcd2 == csr_addr[11:0] ? reg_csr_3282 : _GEN_3281; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3283 = 12'hcd3 == csr_addr[11:0] ? reg_csr_3283 : _GEN_3282; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3284 = 12'hcd4 == csr_addr[11:0] ? reg_csr_3284 : _GEN_3283; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3285 = 12'hcd5 == csr_addr[11:0] ? reg_csr_3285 : _GEN_3284; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3286 = 12'hcd6 == csr_addr[11:0] ? reg_csr_3286 : _GEN_3285; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3287 = 12'hcd7 == csr_addr[11:0] ? reg_csr_3287 : _GEN_3286; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3288 = 12'hcd8 == csr_addr[11:0] ? reg_csr_3288 : _GEN_3287; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3289 = 12'hcd9 == csr_addr[11:0] ? reg_csr_3289 : _GEN_3288; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3290 = 12'hcda == csr_addr[11:0] ? reg_csr_3290 : _GEN_3289; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3291 = 12'hcdb == csr_addr[11:0] ? reg_csr_3291 : _GEN_3290; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3292 = 12'hcdc == csr_addr[11:0] ? reg_csr_3292 : _GEN_3291; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3293 = 12'hcdd == csr_addr[11:0] ? reg_csr_3293 : _GEN_3292; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3294 = 12'hcde == csr_addr[11:0] ? reg_csr_3294 : _GEN_3293; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3295 = 12'hcdf == csr_addr[11:0] ? reg_csr_3295 : _GEN_3294; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3296 = 12'hce0 == csr_addr[11:0] ? reg_csr_3296 : _GEN_3295; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3297 = 12'hce1 == csr_addr[11:0] ? reg_csr_3297 : _GEN_3296; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3298 = 12'hce2 == csr_addr[11:0] ? reg_csr_3298 : _GEN_3297; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3299 = 12'hce3 == csr_addr[11:0] ? reg_csr_3299 : _GEN_3298; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3300 = 12'hce4 == csr_addr[11:0] ? reg_csr_3300 : _GEN_3299; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3301 = 12'hce5 == csr_addr[11:0] ? reg_csr_3301 : _GEN_3300; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3302 = 12'hce6 == csr_addr[11:0] ? reg_csr_3302 : _GEN_3301; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3303 = 12'hce7 == csr_addr[11:0] ? reg_csr_3303 : _GEN_3302; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3304 = 12'hce8 == csr_addr[11:0] ? reg_csr_3304 : _GEN_3303; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3305 = 12'hce9 == csr_addr[11:0] ? reg_csr_3305 : _GEN_3304; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3306 = 12'hcea == csr_addr[11:0] ? reg_csr_3306 : _GEN_3305; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3307 = 12'hceb == csr_addr[11:0] ? reg_csr_3307 : _GEN_3306; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3308 = 12'hcec == csr_addr[11:0] ? reg_csr_3308 : _GEN_3307; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3309 = 12'hced == csr_addr[11:0] ? reg_csr_3309 : _GEN_3308; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3310 = 12'hcee == csr_addr[11:0] ? reg_csr_3310 : _GEN_3309; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3311 = 12'hcef == csr_addr[11:0] ? reg_csr_3311 : _GEN_3310; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3312 = 12'hcf0 == csr_addr[11:0] ? reg_csr_3312 : _GEN_3311; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3313 = 12'hcf1 == csr_addr[11:0] ? reg_csr_3313 : _GEN_3312; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3314 = 12'hcf2 == csr_addr[11:0] ? reg_csr_3314 : _GEN_3313; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3315 = 12'hcf3 == csr_addr[11:0] ? reg_csr_3315 : _GEN_3314; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3316 = 12'hcf4 == csr_addr[11:0] ? reg_csr_3316 : _GEN_3315; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3317 = 12'hcf5 == csr_addr[11:0] ? reg_csr_3317 : _GEN_3316; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3318 = 12'hcf6 == csr_addr[11:0] ? reg_csr_3318 : _GEN_3317; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3319 = 12'hcf7 == csr_addr[11:0] ? reg_csr_3319 : _GEN_3318; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3320 = 12'hcf8 == csr_addr[11:0] ? reg_csr_3320 : _GEN_3319; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3321 = 12'hcf9 == csr_addr[11:0] ? reg_csr_3321 : _GEN_3320; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3322 = 12'hcfa == csr_addr[11:0] ? reg_csr_3322 : _GEN_3321; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3323 = 12'hcfb == csr_addr[11:0] ? reg_csr_3323 : _GEN_3322; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3324 = 12'hcfc == csr_addr[11:0] ? reg_csr_3324 : _GEN_3323; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3325 = 12'hcfd == csr_addr[11:0] ? reg_csr_3325 : _GEN_3324; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3326 = 12'hcfe == csr_addr[11:0] ? reg_csr_3326 : _GEN_3325; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3327 = 12'hcff == csr_addr[11:0] ? reg_csr_3327 : _GEN_3326; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3328 = 12'hd00 == csr_addr[11:0] ? reg_csr_3328 : _GEN_3327; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3329 = 12'hd01 == csr_addr[11:0] ? reg_csr_3329 : _GEN_3328; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3330 = 12'hd02 == csr_addr[11:0] ? reg_csr_3330 : _GEN_3329; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3331 = 12'hd03 == csr_addr[11:0] ? reg_csr_3331 : _GEN_3330; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3332 = 12'hd04 == csr_addr[11:0] ? reg_csr_3332 : _GEN_3331; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3333 = 12'hd05 == csr_addr[11:0] ? reg_csr_3333 : _GEN_3332; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3334 = 12'hd06 == csr_addr[11:0] ? reg_csr_3334 : _GEN_3333; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3335 = 12'hd07 == csr_addr[11:0] ? reg_csr_3335 : _GEN_3334; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3336 = 12'hd08 == csr_addr[11:0] ? reg_csr_3336 : _GEN_3335; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3337 = 12'hd09 == csr_addr[11:0] ? reg_csr_3337 : _GEN_3336; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3338 = 12'hd0a == csr_addr[11:0] ? reg_csr_3338 : _GEN_3337; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3339 = 12'hd0b == csr_addr[11:0] ? reg_csr_3339 : _GEN_3338; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3340 = 12'hd0c == csr_addr[11:0] ? reg_csr_3340 : _GEN_3339; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3341 = 12'hd0d == csr_addr[11:0] ? reg_csr_3341 : _GEN_3340; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3342 = 12'hd0e == csr_addr[11:0] ? reg_csr_3342 : _GEN_3341; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3343 = 12'hd0f == csr_addr[11:0] ? reg_csr_3343 : _GEN_3342; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3344 = 12'hd10 == csr_addr[11:0] ? reg_csr_3344 : _GEN_3343; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3345 = 12'hd11 == csr_addr[11:0] ? reg_csr_3345 : _GEN_3344; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3346 = 12'hd12 == csr_addr[11:0] ? reg_csr_3346 : _GEN_3345; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3347 = 12'hd13 == csr_addr[11:0] ? reg_csr_3347 : _GEN_3346; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3348 = 12'hd14 == csr_addr[11:0] ? reg_csr_3348 : _GEN_3347; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3349 = 12'hd15 == csr_addr[11:0] ? reg_csr_3349 : _GEN_3348; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3350 = 12'hd16 == csr_addr[11:0] ? reg_csr_3350 : _GEN_3349; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3351 = 12'hd17 == csr_addr[11:0] ? reg_csr_3351 : _GEN_3350; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3352 = 12'hd18 == csr_addr[11:0] ? reg_csr_3352 : _GEN_3351; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3353 = 12'hd19 == csr_addr[11:0] ? reg_csr_3353 : _GEN_3352; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3354 = 12'hd1a == csr_addr[11:0] ? reg_csr_3354 : _GEN_3353; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3355 = 12'hd1b == csr_addr[11:0] ? reg_csr_3355 : _GEN_3354; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3356 = 12'hd1c == csr_addr[11:0] ? reg_csr_3356 : _GEN_3355; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3357 = 12'hd1d == csr_addr[11:0] ? reg_csr_3357 : _GEN_3356; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3358 = 12'hd1e == csr_addr[11:0] ? reg_csr_3358 : _GEN_3357; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3359 = 12'hd1f == csr_addr[11:0] ? reg_csr_3359 : _GEN_3358; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3360 = 12'hd20 == csr_addr[11:0] ? reg_csr_3360 : _GEN_3359; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3361 = 12'hd21 == csr_addr[11:0] ? reg_csr_3361 : _GEN_3360; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3362 = 12'hd22 == csr_addr[11:0] ? reg_csr_3362 : _GEN_3361; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3363 = 12'hd23 == csr_addr[11:0] ? reg_csr_3363 : _GEN_3362; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3364 = 12'hd24 == csr_addr[11:0] ? reg_csr_3364 : _GEN_3363; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3365 = 12'hd25 == csr_addr[11:0] ? reg_csr_3365 : _GEN_3364; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3366 = 12'hd26 == csr_addr[11:0] ? reg_csr_3366 : _GEN_3365; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3367 = 12'hd27 == csr_addr[11:0] ? reg_csr_3367 : _GEN_3366; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3368 = 12'hd28 == csr_addr[11:0] ? reg_csr_3368 : _GEN_3367; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3369 = 12'hd29 == csr_addr[11:0] ? reg_csr_3369 : _GEN_3368; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3370 = 12'hd2a == csr_addr[11:0] ? reg_csr_3370 : _GEN_3369; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3371 = 12'hd2b == csr_addr[11:0] ? reg_csr_3371 : _GEN_3370; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3372 = 12'hd2c == csr_addr[11:0] ? reg_csr_3372 : _GEN_3371; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3373 = 12'hd2d == csr_addr[11:0] ? reg_csr_3373 : _GEN_3372; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3374 = 12'hd2e == csr_addr[11:0] ? reg_csr_3374 : _GEN_3373; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3375 = 12'hd2f == csr_addr[11:0] ? reg_csr_3375 : _GEN_3374; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3376 = 12'hd30 == csr_addr[11:0] ? reg_csr_3376 : _GEN_3375; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3377 = 12'hd31 == csr_addr[11:0] ? reg_csr_3377 : _GEN_3376; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3378 = 12'hd32 == csr_addr[11:0] ? reg_csr_3378 : _GEN_3377; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3379 = 12'hd33 == csr_addr[11:0] ? reg_csr_3379 : _GEN_3378; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3380 = 12'hd34 == csr_addr[11:0] ? reg_csr_3380 : _GEN_3379; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3381 = 12'hd35 == csr_addr[11:0] ? reg_csr_3381 : _GEN_3380; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3382 = 12'hd36 == csr_addr[11:0] ? reg_csr_3382 : _GEN_3381; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3383 = 12'hd37 == csr_addr[11:0] ? reg_csr_3383 : _GEN_3382; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3384 = 12'hd38 == csr_addr[11:0] ? reg_csr_3384 : _GEN_3383; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3385 = 12'hd39 == csr_addr[11:0] ? reg_csr_3385 : _GEN_3384; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3386 = 12'hd3a == csr_addr[11:0] ? reg_csr_3386 : _GEN_3385; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3387 = 12'hd3b == csr_addr[11:0] ? reg_csr_3387 : _GEN_3386; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3388 = 12'hd3c == csr_addr[11:0] ? reg_csr_3388 : _GEN_3387; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3389 = 12'hd3d == csr_addr[11:0] ? reg_csr_3389 : _GEN_3388; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3390 = 12'hd3e == csr_addr[11:0] ? reg_csr_3390 : _GEN_3389; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3391 = 12'hd3f == csr_addr[11:0] ? reg_csr_3391 : _GEN_3390; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3392 = 12'hd40 == csr_addr[11:0] ? reg_csr_3392 : _GEN_3391; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3393 = 12'hd41 == csr_addr[11:0] ? reg_csr_3393 : _GEN_3392; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3394 = 12'hd42 == csr_addr[11:0] ? reg_csr_3394 : _GEN_3393; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3395 = 12'hd43 == csr_addr[11:0] ? reg_csr_3395 : _GEN_3394; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3396 = 12'hd44 == csr_addr[11:0] ? reg_csr_3396 : _GEN_3395; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3397 = 12'hd45 == csr_addr[11:0] ? reg_csr_3397 : _GEN_3396; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3398 = 12'hd46 == csr_addr[11:0] ? reg_csr_3398 : _GEN_3397; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3399 = 12'hd47 == csr_addr[11:0] ? reg_csr_3399 : _GEN_3398; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3400 = 12'hd48 == csr_addr[11:0] ? reg_csr_3400 : _GEN_3399; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3401 = 12'hd49 == csr_addr[11:0] ? reg_csr_3401 : _GEN_3400; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3402 = 12'hd4a == csr_addr[11:0] ? reg_csr_3402 : _GEN_3401; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3403 = 12'hd4b == csr_addr[11:0] ? reg_csr_3403 : _GEN_3402; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3404 = 12'hd4c == csr_addr[11:0] ? reg_csr_3404 : _GEN_3403; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3405 = 12'hd4d == csr_addr[11:0] ? reg_csr_3405 : _GEN_3404; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3406 = 12'hd4e == csr_addr[11:0] ? reg_csr_3406 : _GEN_3405; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3407 = 12'hd4f == csr_addr[11:0] ? reg_csr_3407 : _GEN_3406; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3408 = 12'hd50 == csr_addr[11:0] ? reg_csr_3408 : _GEN_3407; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3409 = 12'hd51 == csr_addr[11:0] ? reg_csr_3409 : _GEN_3408; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3410 = 12'hd52 == csr_addr[11:0] ? reg_csr_3410 : _GEN_3409; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3411 = 12'hd53 == csr_addr[11:0] ? reg_csr_3411 : _GEN_3410; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3412 = 12'hd54 == csr_addr[11:0] ? reg_csr_3412 : _GEN_3411; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3413 = 12'hd55 == csr_addr[11:0] ? reg_csr_3413 : _GEN_3412; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3414 = 12'hd56 == csr_addr[11:0] ? reg_csr_3414 : _GEN_3413; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3415 = 12'hd57 == csr_addr[11:0] ? reg_csr_3415 : _GEN_3414; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3416 = 12'hd58 == csr_addr[11:0] ? reg_csr_3416 : _GEN_3415; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3417 = 12'hd59 == csr_addr[11:0] ? reg_csr_3417 : _GEN_3416; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3418 = 12'hd5a == csr_addr[11:0] ? reg_csr_3418 : _GEN_3417; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3419 = 12'hd5b == csr_addr[11:0] ? reg_csr_3419 : _GEN_3418; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3420 = 12'hd5c == csr_addr[11:0] ? reg_csr_3420 : _GEN_3419; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3421 = 12'hd5d == csr_addr[11:0] ? reg_csr_3421 : _GEN_3420; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3422 = 12'hd5e == csr_addr[11:0] ? reg_csr_3422 : _GEN_3421; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3423 = 12'hd5f == csr_addr[11:0] ? reg_csr_3423 : _GEN_3422; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3424 = 12'hd60 == csr_addr[11:0] ? reg_csr_3424 : _GEN_3423; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3425 = 12'hd61 == csr_addr[11:0] ? reg_csr_3425 : _GEN_3424; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3426 = 12'hd62 == csr_addr[11:0] ? reg_csr_3426 : _GEN_3425; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3427 = 12'hd63 == csr_addr[11:0] ? reg_csr_3427 : _GEN_3426; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3428 = 12'hd64 == csr_addr[11:0] ? reg_csr_3428 : _GEN_3427; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3429 = 12'hd65 == csr_addr[11:0] ? reg_csr_3429 : _GEN_3428; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3430 = 12'hd66 == csr_addr[11:0] ? reg_csr_3430 : _GEN_3429; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3431 = 12'hd67 == csr_addr[11:0] ? reg_csr_3431 : _GEN_3430; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3432 = 12'hd68 == csr_addr[11:0] ? reg_csr_3432 : _GEN_3431; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3433 = 12'hd69 == csr_addr[11:0] ? reg_csr_3433 : _GEN_3432; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3434 = 12'hd6a == csr_addr[11:0] ? reg_csr_3434 : _GEN_3433; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3435 = 12'hd6b == csr_addr[11:0] ? reg_csr_3435 : _GEN_3434; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3436 = 12'hd6c == csr_addr[11:0] ? reg_csr_3436 : _GEN_3435; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3437 = 12'hd6d == csr_addr[11:0] ? reg_csr_3437 : _GEN_3436; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3438 = 12'hd6e == csr_addr[11:0] ? reg_csr_3438 : _GEN_3437; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3439 = 12'hd6f == csr_addr[11:0] ? reg_csr_3439 : _GEN_3438; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3440 = 12'hd70 == csr_addr[11:0] ? reg_csr_3440 : _GEN_3439; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3441 = 12'hd71 == csr_addr[11:0] ? reg_csr_3441 : _GEN_3440; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3442 = 12'hd72 == csr_addr[11:0] ? reg_csr_3442 : _GEN_3441; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3443 = 12'hd73 == csr_addr[11:0] ? reg_csr_3443 : _GEN_3442; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3444 = 12'hd74 == csr_addr[11:0] ? reg_csr_3444 : _GEN_3443; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3445 = 12'hd75 == csr_addr[11:0] ? reg_csr_3445 : _GEN_3444; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3446 = 12'hd76 == csr_addr[11:0] ? reg_csr_3446 : _GEN_3445; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3447 = 12'hd77 == csr_addr[11:0] ? reg_csr_3447 : _GEN_3446; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3448 = 12'hd78 == csr_addr[11:0] ? reg_csr_3448 : _GEN_3447; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3449 = 12'hd79 == csr_addr[11:0] ? reg_csr_3449 : _GEN_3448; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3450 = 12'hd7a == csr_addr[11:0] ? reg_csr_3450 : _GEN_3449; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3451 = 12'hd7b == csr_addr[11:0] ? reg_csr_3451 : _GEN_3450; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3452 = 12'hd7c == csr_addr[11:0] ? reg_csr_3452 : _GEN_3451; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3453 = 12'hd7d == csr_addr[11:0] ? reg_csr_3453 : _GEN_3452; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3454 = 12'hd7e == csr_addr[11:0] ? reg_csr_3454 : _GEN_3453; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3455 = 12'hd7f == csr_addr[11:0] ? reg_csr_3455 : _GEN_3454; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3456 = 12'hd80 == csr_addr[11:0] ? reg_csr_3456 : _GEN_3455; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3457 = 12'hd81 == csr_addr[11:0] ? reg_csr_3457 : _GEN_3456; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3458 = 12'hd82 == csr_addr[11:0] ? reg_csr_3458 : _GEN_3457; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3459 = 12'hd83 == csr_addr[11:0] ? reg_csr_3459 : _GEN_3458; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3460 = 12'hd84 == csr_addr[11:0] ? reg_csr_3460 : _GEN_3459; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3461 = 12'hd85 == csr_addr[11:0] ? reg_csr_3461 : _GEN_3460; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3462 = 12'hd86 == csr_addr[11:0] ? reg_csr_3462 : _GEN_3461; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3463 = 12'hd87 == csr_addr[11:0] ? reg_csr_3463 : _GEN_3462; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3464 = 12'hd88 == csr_addr[11:0] ? reg_csr_3464 : _GEN_3463; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3465 = 12'hd89 == csr_addr[11:0] ? reg_csr_3465 : _GEN_3464; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3466 = 12'hd8a == csr_addr[11:0] ? reg_csr_3466 : _GEN_3465; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3467 = 12'hd8b == csr_addr[11:0] ? reg_csr_3467 : _GEN_3466; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3468 = 12'hd8c == csr_addr[11:0] ? reg_csr_3468 : _GEN_3467; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3469 = 12'hd8d == csr_addr[11:0] ? reg_csr_3469 : _GEN_3468; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3470 = 12'hd8e == csr_addr[11:0] ? reg_csr_3470 : _GEN_3469; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3471 = 12'hd8f == csr_addr[11:0] ? reg_csr_3471 : _GEN_3470; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3472 = 12'hd90 == csr_addr[11:0] ? reg_csr_3472 : _GEN_3471; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3473 = 12'hd91 == csr_addr[11:0] ? reg_csr_3473 : _GEN_3472; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3474 = 12'hd92 == csr_addr[11:0] ? reg_csr_3474 : _GEN_3473; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3475 = 12'hd93 == csr_addr[11:0] ? reg_csr_3475 : _GEN_3474; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3476 = 12'hd94 == csr_addr[11:0] ? reg_csr_3476 : _GEN_3475; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3477 = 12'hd95 == csr_addr[11:0] ? reg_csr_3477 : _GEN_3476; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3478 = 12'hd96 == csr_addr[11:0] ? reg_csr_3478 : _GEN_3477; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3479 = 12'hd97 == csr_addr[11:0] ? reg_csr_3479 : _GEN_3478; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3480 = 12'hd98 == csr_addr[11:0] ? reg_csr_3480 : _GEN_3479; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3481 = 12'hd99 == csr_addr[11:0] ? reg_csr_3481 : _GEN_3480; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3482 = 12'hd9a == csr_addr[11:0] ? reg_csr_3482 : _GEN_3481; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3483 = 12'hd9b == csr_addr[11:0] ? reg_csr_3483 : _GEN_3482; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3484 = 12'hd9c == csr_addr[11:0] ? reg_csr_3484 : _GEN_3483; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3485 = 12'hd9d == csr_addr[11:0] ? reg_csr_3485 : _GEN_3484; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3486 = 12'hd9e == csr_addr[11:0] ? reg_csr_3486 : _GEN_3485; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3487 = 12'hd9f == csr_addr[11:0] ? reg_csr_3487 : _GEN_3486; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3488 = 12'hda0 == csr_addr[11:0] ? reg_csr_3488 : _GEN_3487; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3489 = 12'hda1 == csr_addr[11:0] ? reg_csr_3489 : _GEN_3488; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3490 = 12'hda2 == csr_addr[11:0] ? reg_csr_3490 : _GEN_3489; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3491 = 12'hda3 == csr_addr[11:0] ? reg_csr_3491 : _GEN_3490; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3492 = 12'hda4 == csr_addr[11:0] ? reg_csr_3492 : _GEN_3491; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3493 = 12'hda5 == csr_addr[11:0] ? reg_csr_3493 : _GEN_3492; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3494 = 12'hda6 == csr_addr[11:0] ? reg_csr_3494 : _GEN_3493; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3495 = 12'hda7 == csr_addr[11:0] ? reg_csr_3495 : _GEN_3494; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3496 = 12'hda8 == csr_addr[11:0] ? reg_csr_3496 : _GEN_3495; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3497 = 12'hda9 == csr_addr[11:0] ? reg_csr_3497 : _GEN_3496; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3498 = 12'hdaa == csr_addr[11:0] ? reg_csr_3498 : _GEN_3497; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3499 = 12'hdab == csr_addr[11:0] ? reg_csr_3499 : _GEN_3498; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3500 = 12'hdac == csr_addr[11:0] ? reg_csr_3500 : _GEN_3499; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3501 = 12'hdad == csr_addr[11:0] ? reg_csr_3501 : _GEN_3500; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3502 = 12'hdae == csr_addr[11:0] ? reg_csr_3502 : _GEN_3501; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3503 = 12'hdaf == csr_addr[11:0] ? reg_csr_3503 : _GEN_3502; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3504 = 12'hdb0 == csr_addr[11:0] ? reg_csr_3504 : _GEN_3503; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3505 = 12'hdb1 == csr_addr[11:0] ? reg_csr_3505 : _GEN_3504; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3506 = 12'hdb2 == csr_addr[11:0] ? reg_csr_3506 : _GEN_3505; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3507 = 12'hdb3 == csr_addr[11:0] ? reg_csr_3507 : _GEN_3506; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3508 = 12'hdb4 == csr_addr[11:0] ? reg_csr_3508 : _GEN_3507; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3509 = 12'hdb5 == csr_addr[11:0] ? reg_csr_3509 : _GEN_3508; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3510 = 12'hdb6 == csr_addr[11:0] ? reg_csr_3510 : _GEN_3509; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3511 = 12'hdb7 == csr_addr[11:0] ? reg_csr_3511 : _GEN_3510; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3512 = 12'hdb8 == csr_addr[11:0] ? reg_csr_3512 : _GEN_3511; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3513 = 12'hdb9 == csr_addr[11:0] ? reg_csr_3513 : _GEN_3512; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3514 = 12'hdba == csr_addr[11:0] ? reg_csr_3514 : _GEN_3513; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3515 = 12'hdbb == csr_addr[11:0] ? reg_csr_3515 : _GEN_3514; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3516 = 12'hdbc == csr_addr[11:0] ? reg_csr_3516 : _GEN_3515; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3517 = 12'hdbd == csr_addr[11:0] ? reg_csr_3517 : _GEN_3516; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3518 = 12'hdbe == csr_addr[11:0] ? reg_csr_3518 : _GEN_3517; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3519 = 12'hdbf == csr_addr[11:0] ? reg_csr_3519 : _GEN_3518; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3520 = 12'hdc0 == csr_addr[11:0] ? reg_csr_3520 : _GEN_3519; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3521 = 12'hdc1 == csr_addr[11:0] ? reg_csr_3521 : _GEN_3520; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3522 = 12'hdc2 == csr_addr[11:0] ? reg_csr_3522 : _GEN_3521; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3523 = 12'hdc3 == csr_addr[11:0] ? reg_csr_3523 : _GEN_3522; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3524 = 12'hdc4 == csr_addr[11:0] ? reg_csr_3524 : _GEN_3523; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3525 = 12'hdc5 == csr_addr[11:0] ? reg_csr_3525 : _GEN_3524; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3526 = 12'hdc6 == csr_addr[11:0] ? reg_csr_3526 : _GEN_3525; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3527 = 12'hdc7 == csr_addr[11:0] ? reg_csr_3527 : _GEN_3526; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3528 = 12'hdc8 == csr_addr[11:0] ? reg_csr_3528 : _GEN_3527; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3529 = 12'hdc9 == csr_addr[11:0] ? reg_csr_3529 : _GEN_3528; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3530 = 12'hdca == csr_addr[11:0] ? reg_csr_3530 : _GEN_3529; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3531 = 12'hdcb == csr_addr[11:0] ? reg_csr_3531 : _GEN_3530; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3532 = 12'hdcc == csr_addr[11:0] ? reg_csr_3532 : _GEN_3531; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3533 = 12'hdcd == csr_addr[11:0] ? reg_csr_3533 : _GEN_3532; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3534 = 12'hdce == csr_addr[11:0] ? reg_csr_3534 : _GEN_3533; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3535 = 12'hdcf == csr_addr[11:0] ? reg_csr_3535 : _GEN_3534; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3536 = 12'hdd0 == csr_addr[11:0] ? reg_csr_3536 : _GEN_3535; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3537 = 12'hdd1 == csr_addr[11:0] ? reg_csr_3537 : _GEN_3536; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3538 = 12'hdd2 == csr_addr[11:0] ? reg_csr_3538 : _GEN_3537; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3539 = 12'hdd3 == csr_addr[11:0] ? reg_csr_3539 : _GEN_3538; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3540 = 12'hdd4 == csr_addr[11:0] ? reg_csr_3540 : _GEN_3539; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3541 = 12'hdd5 == csr_addr[11:0] ? reg_csr_3541 : _GEN_3540; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3542 = 12'hdd6 == csr_addr[11:0] ? reg_csr_3542 : _GEN_3541; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3543 = 12'hdd7 == csr_addr[11:0] ? reg_csr_3543 : _GEN_3542; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3544 = 12'hdd8 == csr_addr[11:0] ? reg_csr_3544 : _GEN_3543; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3545 = 12'hdd9 == csr_addr[11:0] ? reg_csr_3545 : _GEN_3544; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3546 = 12'hdda == csr_addr[11:0] ? reg_csr_3546 : _GEN_3545; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3547 = 12'hddb == csr_addr[11:0] ? reg_csr_3547 : _GEN_3546; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3548 = 12'hddc == csr_addr[11:0] ? reg_csr_3548 : _GEN_3547; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3549 = 12'hddd == csr_addr[11:0] ? reg_csr_3549 : _GEN_3548; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3550 = 12'hdde == csr_addr[11:0] ? reg_csr_3550 : _GEN_3549; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3551 = 12'hddf == csr_addr[11:0] ? reg_csr_3551 : _GEN_3550; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3552 = 12'hde0 == csr_addr[11:0] ? reg_csr_3552 : _GEN_3551; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3553 = 12'hde1 == csr_addr[11:0] ? reg_csr_3553 : _GEN_3552; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3554 = 12'hde2 == csr_addr[11:0] ? reg_csr_3554 : _GEN_3553; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3555 = 12'hde3 == csr_addr[11:0] ? reg_csr_3555 : _GEN_3554; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3556 = 12'hde4 == csr_addr[11:0] ? reg_csr_3556 : _GEN_3555; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3557 = 12'hde5 == csr_addr[11:0] ? reg_csr_3557 : _GEN_3556; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3558 = 12'hde6 == csr_addr[11:0] ? reg_csr_3558 : _GEN_3557; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3559 = 12'hde7 == csr_addr[11:0] ? reg_csr_3559 : _GEN_3558; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3560 = 12'hde8 == csr_addr[11:0] ? reg_csr_3560 : _GEN_3559; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3561 = 12'hde9 == csr_addr[11:0] ? reg_csr_3561 : _GEN_3560; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3562 = 12'hdea == csr_addr[11:0] ? reg_csr_3562 : _GEN_3561; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3563 = 12'hdeb == csr_addr[11:0] ? reg_csr_3563 : _GEN_3562; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3564 = 12'hdec == csr_addr[11:0] ? reg_csr_3564 : _GEN_3563; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3565 = 12'hded == csr_addr[11:0] ? reg_csr_3565 : _GEN_3564; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3566 = 12'hdee == csr_addr[11:0] ? reg_csr_3566 : _GEN_3565; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3567 = 12'hdef == csr_addr[11:0] ? reg_csr_3567 : _GEN_3566; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3568 = 12'hdf0 == csr_addr[11:0] ? reg_csr_3568 : _GEN_3567; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3569 = 12'hdf1 == csr_addr[11:0] ? reg_csr_3569 : _GEN_3568; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3570 = 12'hdf2 == csr_addr[11:0] ? reg_csr_3570 : _GEN_3569; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3571 = 12'hdf3 == csr_addr[11:0] ? reg_csr_3571 : _GEN_3570; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3572 = 12'hdf4 == csr_addr[11:0] ? reg_csr_3572 : _GEN_3571; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3573 = 12'hdf5 == csr_addr[11:0] ? reg_csr_3573 : _GEN_3572; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3574 = 12'hdf6 == csr_addr[11:0] ? reg_csr_3574 : _GEN_3573; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3575 = 12'hdf7 == csr_addr[11:0] ? reg_csr_3575 : _GEN_3574; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3576 = 12'hdf8 == csr_addr[11:0] ? reg_csr_3576 : _GEN_3575; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3577 = 12'hdf9 == csr_addr[11:0] ? reg_csr_3577 : _GEN_3576; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3578 = 12'hdfa == csr_addr[11:0] ? reg_csr_3578 : _GEN_3577; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3579 = 12'hdfb == csr_addr[11:0] ? reg_csr_3579 : _GEN_3578; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3580 = 12'hdfc == csr_addr[11:0] ? reg_csr_3580 : _GEN_3579; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3581 = 12'hdfd == csr_addr[11:0] ? reg_csr_3581 : _GEN_3580; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3582 = 12'hdfe == csr_addr[11:0] ? reg_csr_3582 : _GEN_3581; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3583 = 12'hdff == csr_addr[11:0] ? reg_csr_3583 : _GEN_3582; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3584 = 12'he00 == csr_addr[11:0] ? reg_csr_3584 : _GEN_3583; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3585 = 12'he01 == csr_addr[11:0] ? reg_csr_3585 : _GEN_3584; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3586 = 12'he02 == csr_addr[11:0] ? reg_csr_3586 : _GEN_3585; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3587 = 12'he03 == csr_addr[11:0] ? reg_csr_3587 : _GEN_3586; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3588 = 12'he04 == csr_addr[11:0] ? reg_csr_3588 : _GEN_3587; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3589 = 12'he05 == csr_addr[11:0] ? reg_csr_3589 : _GEN_3588; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3590 = 12'he06 == csr_addr[11:0] ? reg_csr_3590 : _GEN_3589; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3591 = 12'he07 == csr_addr[11:0] ? reg_csr_3591 : _GEN_3590; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3592 = 12'he08 == csr_addr[11:0] ? reg_csr_3592 : _GEN_3591; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3593 = 12'he09 == csr_addr[11:0] ? reg_csr_3593 : _GEN_3592; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3594 = 12'he0a == csr_addr[11:0] ? reg_csr_3594 : _GEN_3593; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3595 = 12'he0b == csr_addr[11:0] ? reg_csr_3595 : _GEN_3594; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3596 = 12'he0c == csr_addr[11:0] ? reg_csr_3596 : _GEN_3595; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3597 = 12'he0d == csr_addr[11:0] ? reg_csr_3597 : _GEN_3596; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3598 = 12'he0e == csr_addr[11:0] ? reg_csr_3598 : _GEN_3597; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3599 = 12'he0f == csr_addr[11:0] ? reg_csr_3599 : _GEN_3598; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3600 = 12'he10 == csr_addr[11:0] ? reg_csr_3600 : _GEN_3599; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3601 = 12'he11 == csr_addr[11:0] ? reg_csr_3601 : _GEN_3600; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3602 = 12'he12 == csr_addr[11:0] ? reg_csr_3602 : _GEN_3601; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3603 = 12'he13 == csr_addr[11:0] ? reg_csr_3603 : _GEN_3602; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3604 = 12'he14 == csr_addr[11:0] ? reg_csr_3604 : _GEN_3603; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3605 = 12'he15 == csr_addr[11:0] ? reg_csr_3605 : _GEN_3604; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3606 = 12'he16 == csr_addr[11:0] ? reg_csr_3606 : _GEN_3605; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3607 = 12'he17 == csr_addr[11:0] ? reg_csr_3607 : _GEN_3606; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3608 = 12'he18 == csr_addr[11:0] ? reg_csr_3608 : _GEN_3607; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3609 = 12'he19 == csr_addr[11:0] ? reg_csr_3609 : _GEN_3608; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3610 = 12'he1a == csr_addr[11:0] ? reg_csr_3610 : _GEN_3609; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3611 = 12'he1b == csr_addr[11:0] ? reg_csr_3611 : _GEN_3610; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3612 = 12'he1c == csr_addr[11:0] ? reg_csr_3612 : _GEN_3611; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3613 = 12'he1d == csr_addr[11:0] ? reg_csr_3613 : _GEN_3612; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3614 = 12'he1e == csr_addr[11:0] ? reg_csr_3614 : _GEN_3613; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3615 = 12'he1f == csr_addr[11:0] ? reg_csr_3615 : _GEN_3614; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3616 = 12'he20 == csr_addr[11:0] ? reg_csr_3616 : _GEN_3615; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3617 = 12'he21 == csr_addr[11:0] ? reg_csr_3617 : _GEN_3616; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3618 = 12'he22 == csr_addr[11:0] ? reg_csr_3618 : _GEN_3617; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3619 = 12'he23 == csr_addr[11:0] ? reg_csr_3619 : _GEN_3618; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3620 = 12'he24 == csr_addr[11:0] ? reg_csr_3620 : _GEN_3619; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3621 = 12'he25 == csr_addr[11:0] ? reg_csr_3621 : _GEN_3620; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3622 = 12'he26 == csr_addr[11:0] ? reg_csr_3622 : _GEN_3621; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3623 = 12'he27 == csr_addr[11:0] ? reg_csr_3623 : _GEN_3622; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3624 = 12'he28 == csr_addr[11:0] ? reg_csr_3624 : _GEN_3623; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3625 = 12'he29 == csr_addr[11:0] ? reg_csr_3625 : _GEN_3624; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3626 = 12'he2a == csr_addr[11:0] ? reg_csr_3626 : _GEN_3625; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3627 = 12'he2b == csr_addr[11:0] ? reg_csr_3627 : _GEN_3626; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3628 = 12'he2c == csr_addr[11:0] ? reg_csr_3628 : _GEN_3627; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3629 = 12'he2d == csr_addr[11:0] ? reg_csr_3629 : _GEN_3628; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3630 = 12'he2e == csr_addr[11:0] ? reg_csr_3630 : _GEN_3629; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3631 = 12'he2f == csr_addr[11:0] ? reg_csr_3631 : _GEN_3630; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3632 = 12'he30 == csr_addr[11:0] ? reg_csr_3632 : _GEN_3631; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3633 = 12'he31 == csr_addr[11:0] ? reg_csr_3633 : _GEN_3632; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3634 = 12'he32 == csr_addr[11:0] ? reg_csr_3634 : _GEN_3633; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3635 = 12'he33 == csr_addr[11:0] ? reg_csr_3635 : _GEN_3634; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3636 = 12'he34 == csr_addr[11:0] ? reg_csr_3636 : _GEN_3635; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3637 = 12'he35 == csr_addr[11:0] ? reg_csr_3637 : _GEN_3636; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3638 = 12'he36 == csr_addr[11:0] ? reg_csr_3638 : _GEN_3637; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3639 = 12'he37 == csr_addr[11:0] ? reg_csr_3639 : _GEN_3638; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3640 = 12'he38 == csr_addr[11:0] ? reg_csr_3640 : _GEN_3639; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3641 = 12'he39 == csr_addr[11:0] ? reg_csr_3641 : _GEN_3640; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3642 = 12'he3a == csr_addr[11:0] ? reg_csr_3642 : _GEN_3641; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3643 = 12'he3b == csr_addr[11:0] ? reg_csr_3643 : _GEN_3642; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3644 = 12'he3c == csr_addr[11:0] ? reg_csr_3644 : _GEN_3643; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3645 = 12'he3d == csr_addr[11:0] ? reg_csr_3645 : _GEN_3644; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3646 = 12'he3e == csr_addr[11:0] ? reg_csr_3646 : _GEN_3645; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3647 = 12'he3f == csr_addr[11:0] ? reg_csr_3647 : _GEN_3646; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3648 = 12'he40 == csr_addr[11:0] ? reg_csr_3648 : _GEN_3647; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3649 = 12'he41 == csr_addr[11:0] ? reg_csr_3649 : _GEN_3648; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3650 = 12'he42 == csr_addr[11:0] ? reg_csr_3650 : _GEN_3649; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3651 = 12'he43 == csr_addr[11:0] ? reg_csr_3651 : _GEN_3650; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3652 = 12'he44 == csr_addr[11:0] ? reg_csr_3652 : _GEN_3651; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3653 = 12'he45 == csr_addr[11:0] ? reg_csr_3653 : _GEN_3652; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3654 = 12'he46 == csr_addr[11:0] ? reg_csr_3654 : _GEN_3653; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3655 = 12'he47 == csr_addr[11:0] ? reg_csr_3655 : _GEN_3654; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3656 = 12'he48 == csr_addr[11:0] ? reg_csr_3656 : _GEN_3655; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3657 = 12'he49 == csr_addr[11:0] ? reg_csr_3657 : _GEN_3656; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3658 = 12'he4a == csr_addr[11:0] ? reg_csr_3658 : _GEN_3657; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3659 = 12'he4b == csr_addr[11:0] ? reg_csr_3659 : _GEN_3658; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3660 = 12'he4c == csr_addr[11:0] ? reg_csr_3660 : _GEN_3659; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3661 = 12'he4d == csr_addr[11:0] ? reg_csr_3661 : _GEN_3660; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3662 = 12'he4e == csr_addr[11:0] ? reg_csr_3662 : _GEN_3661; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3663 = 12'he4f == csr_addr[11:0] ? reg_csr_3663 : _GEN_3662; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3664 = 12'he50 == csr_addr[11:0] ? reg_csr_3664 : _GEN_3663; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3665 = 12'he51 == csr_addr[11:0] ? reg_csr_3665 : _GEN_3664; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3666 = 12'he52 == csr_addr[11:0] ? reg_csr_3666 : _GEN_3665; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3667 = 12'he53 == csr_addr[11:0] ? reg_csr_3667 : _GEN_3666; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3668 = 12'he54 == csr_addr[11:0] ? reg_csr_3668 : _GEN_3667; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3669 = 12'he55 == csr_addr[11:0] ? reg_csr_3669 : _GEN_3668; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3670 = 12'he56 == csr_addr[11:0] ? reg_csr_3670 : _GEN_3669; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3671 = 12'he57 == csr_addr[11:0] ? reg_csr_3671 : _GEN_3670; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3672 = 12'he58 == csr_addr[11:0] ? reg_csr_3672 : _GEN_3671; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3673 = 12'he59 == csr_addr[11:0] ? reg_csr_3673 : _GEN_3672; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3674 = 12'he5a == csr_addr[11:0] ? reg_csr_3674 : _GEN_3673; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3675 = 12'he5b == csr_addr[11:0] ? reg_csr_3675 : _GEN_3674; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3676 = 12'he5c == csr_addr[11:0] ? reg_csr_3676 : _GEN_3675; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3677 = 12'he5d == csr_addr[11:0] ? reg_csr_3677 : _GEN_3676; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3678 = 12'he5e == csr_addr[11:0] ? reg_csr_3678 : _GEN_3677; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3679 = 12'he5f == csr_addr[11:0] ? reg_csr_3679 : _GEN_3678; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3680 = 12'he60 == csr_addr[11:0] ? reg_csr_3680 : _GEN_3679; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3681 = 12'he61 == csr_addr[11:0] ? reg_csr_3681 : _GEN_3680; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3682 = 12'he62 == csr_addr[11:0] ? reg_csr_3682 : _GEN_3681; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3683 = 12'he63 == csr_addr[11:0] ? reg_csr_3683 : _GEN_3682; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3684 = 12'he64 == csr_addr[11:0] ? reg_csr_3684 : _GEN_3683; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3685 = 12'he65 == csr_addr[11:0] ? reg_csr_3685 : _GEN_3684; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3686 = 12'he66 == csr_addr[11:0] ? reg_csr_3686 : _GEN_3685; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3687 = 12'he67 == csr_addr[11:0] ? reg_csr_3687 : _GEN_3686; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3688 = 12'he68 == csr_addr[11:0] ? reg_csr_3688 : _GEN_3687; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3689 = 12'he69 == csr_addr[11:0] ? reg_csr_3689 : _GEN_3688; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3690 = 12'he6a == csr_addr[11:0] ? reg_csr_3690 : _GEN_3689; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3691 = 12'he6b == csr_addr[11:0] ? reg_csr_3691 : _GEN_3690; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3692 = 12'he6c == csr_addr[11:0] ? reg_csr_3692 : _GEN_3691; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3693 = 12'he6d == csr_addr[11:0] ? reg_csr_3693 : _GEN_3692; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3694 = 12'he6e == csr_addr[11:0] ? reg_csr_3694 : _GEN_3693; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3695 = 12'he6f == csr_addr[11:0] ? reg_csr_3695 : _GEN_3694; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3696 = 12'he70 == csr_addr[11:0] ? reg_csr_3696 : _GEN_3695; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3697 = 12'he71 == csr_addr[11:0] ? reg_csr_3697 : _GEN_3696; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3698 = 12'he72 == csr_addr[11:0] ? reg_csr_3698 : _GEN_3697; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3699 = 12'he73 == csr_addr[11:0] ? reg_csr_3699 : _GEN_3698; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3700 = 12'he74 == csr_addr[11:0] ? reg_csr_3700 : _GEN_3699; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3701 = 12'he75 == csr_addr[11:0] ? reg_csr_3701 : _GEN_3700; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3702 = 12'he76 == csr_addr[11:0] ? reg_csr_3702 : _GEN_3701; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3703 = 12'he77 == csr_addr[11:0] ? reg_csr_3703 : _GEN_3702; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3704 = 12'he78 == csr_addr[11:0] ? reg_csr_3704 : _GEN_3703; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3705 = 12'he79 == csr_addr[11:0] ? reg_csr_3705 : _GEN_3704; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3706 = 12'he7a == csr_addr[11:0] ? reg_csr_3706 : _GEN_3705; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3707 = 12'he7b == csr_addr[11:0] ? reg_csr_3707 : _GEN_3706; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3708 = 12'he7c == csr_addr[11:0] ? reg_csr_3708 : _GEN_3707; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3709 = 12'he7d == csr_addr[11:0] ? reg_csr_3709 : _GEN_3708; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3710 = 12'he7e == csr_addr[11:0] ? reg_csr_3710 : _GEN_3709; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3711 = 12'he7f == csr_addr[11:0] ? reg_csr_3711 : _GEN_3710; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3712 = 12'he80 == csr_addr[11:0] ? reg_csr_3712 : _GEN_3711; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3713 = 12'he81 == csr_addr[11:0] ? reg_csr_3713 : _GEN_3712; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3714 = 12'he82 == csr_addr[11:0] ? reg_csr_3714 : _GEN_3713; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3715 = 12'he83 == csr_addr[11:0] ? reg_csr_3715 : _GEN_3714; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3716 = 12'he84 == csr_addr[11:0] ? reg_csr_3716 : _GEN_3715; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3717 = 12'he85 == csr_addr[11:0] ? reg_csr_3717 : _GEN_3716; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3718 = 12'he86 == csr_addr[11:0] ? reg_csr_3718 : _GEN_3717; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3719 = 12'he87 == csr_addr[11:0] ? reg_csr_3719 : _GEN_3718; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3720 = 12'he88 == csr_addr[11:0] ? reg_csr_3720 : _GEN_3719; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3721 = 12'he89 == csr_addr[11:0] ? reg_csr_3721 : _GEN_3720; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3722 = 12'he8a == csr_addr[11:0] ? reg_csr_3722 : _GEN_3721; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3723 = 12'he8b == csr_addr[11:0] ? reg_csr_3723 : _GEN_3722; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3724 = 12'he8c == csr_addr[11:0] ? reg_csr_3724 : _GEN_3723; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3725 = 12'he8d == csr_addr[11:0] ? reg_csr_3725 : _GEN_3724; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3726 = 12'he8e == csr_addr[11:0] ? reg_csr_3726 : _GEN_3725; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3727 = 12'he8f == csr_addr[11:0] ? reg_csr_3727 : _GEN_3726; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3728 = 12'he90 == csr_addr[11:0] ? reg_csr_3728 : _GEN_3727; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3729 = 12'he91 == csr_addr[11:0] ? reg_csr_3729 : _GEN_3728; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3730 = 12'he92 == csr_addr[11:0] ? reg_csr_3730 : _GEN_3729; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3731 = 12'he93 == csr_addr[11:0] ? reg_csr_3731 : _GEN_3730; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3732 = 12'he94 == csr_addr[11:0] ? reg_csr_3732 : _GEN_3731; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3733 = 12'he95 == csr_addr[11:0] ? reg_csr_3733 : _GEN_3732; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3734 = 12'he96 == csr_addr[11:0] ? reg_csr_3734 : _GEN_3733; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3735 = 12'he97 == csr_addr[11:0] ? reg_csr_3735 : _GEN_3734; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3736 = 12'he98 == csr_addr[11:0] ? reg_csr_3736 : _GEN_3735; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3737 = 12'he99 == csr_addr[11:0] ? reg_csr_3737 : _GEN_3736; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3738 = 12'he9a == csr_addr[11:0] ? reg_csr_3738 : _GEN_3737; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3739 = 12'he9b == csr_addr[11:0] ? reg_csr_3739 : _GEN_3738; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3740 = 12'he9c == csr_addr[11:0] ? reg_csr_3740 : _GEN_3739; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3741 = 12'he9d == csr_addr[11:0] ? reg_csr_3741 : _GEN_3740; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3742 = 12'he9e == csr_addr[11:0] ? reg_csr_3742 : _GEN_3741; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3743 = 12'he9f == csr_addr[11:0] ? reg_csr_3743 : _GEN_3742; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3744 = 12'hea0 == csr_addr[11:0] ? reg_csr_3744 : _GEN_3743; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3745 = 12'hea1 == csr_addr[11:0] ? reg_csr_3745 : _GEN_3744; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3746 = 12'hea2 == csr_addr[11:0] ? reg_csr_3746 : _GEN_3745; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3747 = 12'hea3 == csr_addr[11:0] ? reg_csr_3747 : _GEN_3746; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3748 = 12'hea4 == csr_addr[11:0] ? reg_csr_3748 : _GEN_3747; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3749 = 12'hea5 == csr_addr[11:0] ? reg_csr_3749 : _GEN_3748; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3750 = 12'hea6 == csr_addr[11:0] ? reg_csr_3750 : _GEN_3749; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3751 = 12'hea7 == csr_addr[11:0] ? reg_csr_3751 : _GEN_3750; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3752 = 12'hea8 == csr_addr[11:0] ? reg_csr_3752 : _GEN_3751; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3753 = 12'hea9 == csr_addr[11:0] ? reg_csr_3753 : _GEN_3752; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3754 = 12'heaa == csr_addr[11:0] ? reg_csr_3754 : _GEN_3753; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3755 = 12'heab == csr_addr[11:0] ? reg_csr_3755 : _GEN_3754; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3756 = 12'heac == csr_addr[11:0] ? reg_csr_3756 : _GEN_3755; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3757 = 12'head == csr_addr[11:0] ? reg_csr_3757 : _GEN_3756; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3758 = 12'heae == csr_addr[11:0] ? reg_csr_3758 : _GEN_3757; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3759 = 12'heaf == csr_addr[11:0] ? reg_csr_3759 : _GEN_3758; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3760 = 12'heb0 == csr_addr[11:0] ? reg_csr_3760 : _GEN_3759; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3761 = 12'heb1 == csr_addr[11:0] ? reg_csr_3761 : _GEN_3760; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3762 = 12'heb2 == csr_addr[11:0] ? reg_csr_3762 : _GEN_3761; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3763 = 12'heb3 == csr_addr[11:0] ? reg_csr_3763 : _GEN_3762; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3764 = 12'heb4 == csr_addr[11:0] ? reg_csr_3764 : _GEN_3763; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3765 = 12'heb5 == csr_addr[11:0] ? reg_csr_3765 : _GEN_3764; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3766 = 12'heb6 == csr_addr[11:0] ? reg_csr_3766 : _GEN_3765; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3767 = 12'heb7 == csr_addr[11:0] ? reg_csr_3767 : _GEN_3766; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3768 = 12'heb8 == csr_addr[11:0] ? reg_csr_3768 : _GEN_3767; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3769 = 12'heb9 == csr_addr[11:0] ? reg_csr_3769 : _GEN_3768; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3770 = 12'heba == csr_addr[11:0] ? reg_csr_3770 : _GEN_3769; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3771 = 12'hebb == csr_addr[11:0] ? reg_csr_3771 : _GEN_3770; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3772 = 12'hebc == csr_addr[11:0] ? reg_csr_3772 : _GEN_3771; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3773 = 12'hebd == csr_addr[11:0] ? reg_csr_3773 : _GEN_3772; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3774 = 12'hebe == csr_addr[11:0] ? reg_csr_3774 : _GEN_3773; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3775 = 12'hebf == csr_addr[11:0] ? reg_csr_3775 : _GEN_3774; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3776 = 12'hec0 == csr_addr[11:0] ? reg_csr_3776 : _GEN_3775; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3777 = 12'hec1 == csr_addr[11:0] ? reg_csr_3777 : _GEN_3776; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3778 = 12'hec2 == csr_addr[11:0] ? reg_csr_3778 : _GEN_3777; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3779 = 12'hec3 == csr_addr[11:0] ? reg_csr_3779 : _GEN_3778; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3780 = 12'hec4 == csr_addr[11:0] ? reg_csr_3780 : _GEN_3779; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3781 = 12'hec5 == csr_addr[11:0] ? reg_csr_3781 : _GEN_3780; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3782 = 12'hec6 == csr_addr[11:0] ? reg_csr_3782 : _GEN_3781; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3783 = 12'hec7 == csr_addr[11:0] ? reg_csr_3783 : _GEN_3782; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3784 = 12'hec8 == csr_addr[11:0] ? reg_csr_3784 : _GEN_3783; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3785 = 12'hec9 == csr_addr[11:0] ? reg_csr_3785 : _GEN_3784; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3786 = 12'heca == csr_addr[11:0] ? reg_csr_3786 : _GEN_3785; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3787 = 12'hecb == csr_addr[11:0] ? reg_csr_3787 : _GEN_3786; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3788 = 12'hecc == csr_addr[11:0] ? reg_csr_3788 : _GEN_3787; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3789 = 12'hecd == csr_addr[11:0] ? reg_csr_3789 : _GEN_3788; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3790 = 12'hece == csr_addr[11:0] ? reg_csr_3790 : _GEN_3789; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3791 = 12'hecf == csr_addr[11:0] ? reg_csr_3791 : _GEN_3790; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3792 = 12'hed0 == csr_addr[11:0] ? reg_csr_3792 : _GEN_3791; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3793 = 12'hed1 == csr_addr[11:0] ? reg_csr_3793 : _GEN_3792; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3794 = 12'hed2 == csr_addr[11:0] ? reg_csr_3794 : _GEN_3793; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3795 = 12'hed3 == csr_addr[11:0] ? reg_csr_3795 : _GEN_3794; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3796 = 12'hed4 == csr_addr[11:0] ? reg_csr_3796 : _GEN_3795; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3797 = 12'hed5 == csr_addr[11:0] ? reg_csr_3797 : _GEN_3796; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3798 = 12'hed6 == csr_addr[11:0] ? reg_csr_3798 : _GEN_3797; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3799 = 12'hed7 == csr_addr[11:0] ? reg_csr_3799 : _GEN_3798; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3800 = 12'hed8 == csr_addr[11:0] ? reg_csr_3800 : _GEN_3799; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3801 = 12'hed9 == csr_addr[11:0] ? reg_csr_3801 : _GEN_3800; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3802 = 12'heda == csr_addr[11:0] ? reg_csr_3802 : _GEN_3801; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3803 = 12'hedb == csr_addr[11:0] ? reg_csr_3803 : _GEN_3802; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3804 = 12'hedc == csr_addr[11:0] ? reg_csr_3804 : _GEN_3803; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3805 = 12'hedd == csr_addr[11:0] ? reg_csr_3805 : _GEN_3804; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3806 = 12'hede == csr_addr[11:0] ? reg_csr_3806 : _GEN_3805; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3807 = 12'hedf == csr_addr[11:0] ? reg_csr_3807 : _GEN_3806; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3808 = 12'hee0 == csr_addr[11:0] ? reg_csr_3808 : _GEN_3807; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3809 = 12'hee1 == csr_addr[11:0] ? reg_csr_3809 : _GEN_3808; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3810 = 12'hee2 == csr_addr[11:0] ? reg_csr_3810 : _GEN_3809; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3811 = 12'hee3 == csr_addr[11:0] ? reg_csr_3811 : _GEN_3810; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3812 = 12'hee4 == csr_addr[11:0] ? reg_csr_3812 : _GEN_3811; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3813 = 12'hee5 == csr_addr[11:0] ? reg_csr_3813 : _GEN_3812; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3814 = 12'hee6 == csr_addr[11:0] ? reg_csr_3814 : _GEN_3813; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3815 = 12'hee7 == csr_addr[11:0] ? reg_csr_3815 : _GEN_3814; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3816 = 12'hee8 == csr_addr[11:0] ? reg_csr_3816 : _GEN_3815; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3817 = 12'hee9 == csr_addr[11:0] ? reg_csr_3817 : _GEN_3816; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3818 = 12'heea == csr_addr[11:0] ? reg_csr_3818 : _GEN_3817; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3819 = 12'heeb == csr_addr[11:0] ? reg_csr_3819 : _GEN_3818; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3820 = 12'heec == csr_addr[11:0] ? reg_csr_3820 : _GEN_3819; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3821 = 12'heed == csr_addr[11:0] ? reg_csr_3821 : _GEN_3820; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3822 = 12'heee == csr_addr[11:0] ? reg_csr_3822 : _GEN_3821; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3823 = 12'heef == csr_addr[11:0] ? reg_csr_3823 : _GEN_3822; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3824 = 12'hef0 == csr_addr[11:0] ? reg_csr_3824 : _GEN_3823; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3825 = 12'hef1 == csr_addr[11:0] ? reg_csr_3825 : _GEN_3824; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3826 = 12'hef2 == csr_addr[11:0] ? reg_csr_3826 : _GEN_3825; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3827 = 12'hef3 == csr_addr[11:0] ? reg_csr_3827 : _GEN_3826; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3828 = 12'hef4 == csr_addr[11:0] ? reg_csr_3828 : _GEN_3827; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3829 = 12'hef5 == csr_addr[11:0] ? reg_csr_3829 : _GEN_3828; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3830 = 12'hef6 == csr_addr[11:0] ? reg_csr_3830 : _GEN_3829; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3831 = 12'hef7 == csr_addr[11:0] ? reg_csr_3831 : _GEN_3830; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3832 = 12'hef8 == csr_addr[11:0] ? reg_csr_3832 : _GEN_3831; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3833 = 12'hef9 == csr_addr[11:0] ? reg_csr_3833 : _GEN_3832; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3834 = 12'hefa == csr_addr[11:0] ? reg_csr_3834 : _GEN_3833; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3835 = 12'hefb == csr_addr[11:0] ? reg_csr_3835 : _GEN_3834; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3836 = 12'hefc == csr_addr[11:0] ? reg_csr_3836 : _GEN_3835; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3837 = 12'hefd == csr_addr[11:0] ? reg_csr_3837 : _GEN_3836; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3838 = 12'hefe == csr_addr[11:0] ? reg_csr_3838 : _GEN_3837; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3839 = 12'heff == csr_addr[11:0] ? reg_csr_3839 : _GEN_3838; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3840 = 12'hf00 == csr_addr[11:0] ? reg_csr_3840 : _GEN_3839; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3841 = 12'hf01 == csr_addr[11:0] ? reg_csr_3841 : _GEN_3840; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3842 = 12'hf02 == csr_addr[11:0] ? reg_csr_3842 : _GEN_3841; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3843 = 12'hf03 == csr_addr[11:0] ? reg_csr_3843 : _GEN_3842; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3844 = 12'hf04 == csr_addr[11:0] ? reg_csr_3844 : _GEN_3843; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3845 = 12'hf05 == csr_addr[11:0] ? reg_csr_3845 : _GEN_3844; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3846 = 12'hf06 == csr_addr[11:0] ? reg_csr_3846 : _GEN_3845; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3847 = 12'hf07 == csr_addr[11:0] ? reg_csr_3847 : _GEN_3846; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3848 = 12'hf08 == csr_addr[11:0] ? reg_csr_3848 : _GEN_3847; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3849 = 12'hf09 == csr_addr[11:0] ? reg_csr_3849 : _GEN_3848; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3850 = 12'hf0a == csr_addr[11:0] ? reg_csr_3850 : _GEN_3849; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3851 = 12'hf0b == csr_addr[11:0] ? reg_csr_3851 : _GEN_3850; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3852 = 12'hf0c == csr_addr[11:0] ? reg_csr_3852 : _GEN_3851; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3853 = 12'hf0d == csr_addr[11:0] ? reg_csr_3853 : _GEN_3852; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3854 = 12'hf0e == csr_addr[11:0] ? reg_csr_3854 : _GEN_3853; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3855 = 12'hf0f == csr_addr[11:0] ? reg_csr_3855 : _GEN_3854; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3856 = 12'hf10 == csr_addr[11:0] ? reg_csr_3856 : _GEN_3855; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3857 = 12'hf11 == csr_addr[11:0] ? reg_csr_3857 : _GEN_3856; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3858 = 12'hf12 == csr_addr[11:0] ? reg_csr_3858 : _GEN_3857; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3859 = 12'hf13 == csr_addr[11:0] ? reg_csr_3859 : _GEN_3858; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3860 = 12'hf14 == csr_addr[11:0] ? reg_csr_3860 : _GEN_3859; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3861 = 12'hf15 == csr_addr[11:0] ? reg_csr_3861 : _GEN_3860; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3862 = 12'hf16 == csr_addr[11:0] ? reg_csr_3862 : _GEN_3861; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3863 = 12'hf17 == csr_addr[11:0] ? reg_csr_3863 : _GEN_3862; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3864 = 12'hf18 == csr_addr[11:0] ? reg_csr_3864 : _GEN_3863; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3865 = 12'hf19 == csr_addr[11:0] ? reg_csr_3865 : _GEN_3864; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3866 = 12'hf1a == csr_addr[11:0] ? reg_csr_3866 : _GEN_3865; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3867 = 12'hf1b == csr_addr[11:0] ? reg_csr_3867 : _GEN_3866; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3868 = 12'hf1c == csr_addr[11:0] ? reg_csr_3868 : _GEN_3867; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3869 = 12'hf1d == csr_addr[11:0] ? reg_csr_3869 : _GEN_3868; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3870 = 12'hf1e == csr_addr[11:0] ? reg_csr_3870 : _GEN_3869; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3871 = 12'hf1f == csr_addr[11:0] ? reg_csr_3871 : _GEN_3870; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3872 = 12'hf20 == csr_addr[11:0] ? reg_csr_3872 : _GEN_3871; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3873 = 12'hf21 == csr_addr[11:0] ? reg_csr_3873 : _GEN_3872; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3874 = 12'hf22 == csr_addr[11:0] ? reg_csr_3874 : _GEN_3873; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3875 = 12'hf23 == csr_addr[11:0] ? reg_csr_3875 : _GEN_3874; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3876 = 12'hf24 == csr_addr[11:0] ? reg_csr_3876 : _GEN_3875; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3877 = 12'hf25 == csr_addr[11:0] ? reg_csr_3877 : _GEN_3876; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3878 = 12'hf26 == csr_addr[11:0] ? reg_csr_3878 : _GEN_3877; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3879 = 12'hf27 == csr_addr[11:0] ? reg_csr_3879 : _GEN_3878; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3880 = 12'hf28 == csr_addr[11:0] ? reg_csr_3880 : _GEN_3879; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3881 = 12'hf29 == csr_addr[11:0] ? reg_csr_3881 : _GEN_3880; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3882 = 12'hf2a == csr_addr[11:0] ? reg_csr_3882 : _GEN_3881; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3883 = 12'hf2b == csr_addr[11:0] ? reg_csr_3883 : _GEN_3882; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3884 = 12'hf2c == csr_addr[11:0] ? reg_csr_3884 : _GEN_3883; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3885 = 12'hf2d == csr_addr[11:0] ? reg_csr_3885 : _GEN_3884; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3886 = 12'hf2e == csr_addr[11:0] ? reg_csr_3886 : _GEN_3885; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3887 = 12'hf2f == csr_addr[11:0] ? reg_csr_3887 : _GEN_3886; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3888 = 12'hf30 == csr_addr[11:0] ? reg_csr_3888 : _GEN_3887; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3889 = 12'hf31 == csr_addr[11:0] ? reg_csr_3889 : _GEN_3888; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3890 = 12'hf32 == csr_addr[11:0] ? reg_csr_3890 : _GEN_3889; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3891 = 12'hf33 == csr_addr[11:0] ? reg_csr_3891 : _GEN_3890; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3892 = 12'hf34 == csr_addr[11:0] ? reg_csr_3892 : _GEN_3891; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3893 = 12'hf35 == csr_addr[11:0] ? reg_csr_3893 : _GEN_3892; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3894 = 12'hf36 == csr_addr[11:0] ? reg_csr_3894 : _GEN_3893; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3895 = 12'hf37 == csr_addr[11:0] ? reg_csr_3895 : _GEN_3894; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3896 = 12'hf38 == csr_addr[11:0] ? reg_csr_3896 : _GEN_3895; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3897 = 12'hf39 == csr_addr[11:0] ? reg_csr_3897 : _GEN_3896; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3898 = 12'hf3a == csr_addr[11:0] ? reg_csr_3898 : _GEN_3897; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3899 = 12'hf3b == csr_addr[11:0] ? reg_csr_3899 : _GEN_3898; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3900 = 12'hf3c == csr_addr[11:0] ? reg_csr_3900 : _GEN_3899; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3901 = 12'hf3d == csr_addr[11:0] ? reg_csr_3901 : _GEN_3900; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3902 = 12'hf3e == csr_addr[11:0] ? reg_csr_3902 : _GEN_3901; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3903 = 12'hf3f == csr_addr[11:0] ? reg_csr_3903 : _GEN_3902; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3904 = 12'hf40 == csr_addr[11:0] ? reg_csr_3904 : _GEN_3903; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3905 = 12'hf41 == csr_addr[11:0] ? reg_csr_3905 : _GEN_3904; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3906 = 12'hf42 == csr_addr[11:0] ? reg_csr_3906 : _GEN_3905; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3907 = 12'hf43 == csr_addr[11:0] ? reg_csr_3907 : _GEN_3906; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3908 = 12'hf44 == csr_addr[11:0] ? reg_csr_3908 : _GEN_3907; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3909 = 12'hf45 == csr_addr[11:0] ? reg_csr_3909 : _GEN_3908; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3910 = 12'hf46 == csr_addr[11:0] ? reg_csr_3910 : _GEN_3909; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3911 = 12'hf47 == csr_addr[11:0] ? reg_csr_3911 : _GEN_3910; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3912 = 12'hf48 == csr_addr[11:0] ? reg_csr_3912 : _GEN_3911; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3913 = 12'hf49 == csr_addr[11:0] ? reg_csr_3913 : _GEN_3912; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3914 = 12'hf4a == csr_addr[11:0] ? reg_csr_3914 : _GEN_3913; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3915 = 12'hf4b == csr_addr[11:0] ? reg_csr_3915 : _GEN_3914; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3916 = 12'hf4c == csr_addr[11:0] ? reg_csr_3916 : _GEN_3915; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3917 = 12'hf4d == csr_addr[11:0] ? reg_csr_3917 : _GEN_3916; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3918 = 12'hf4e == csr_addr[11:0] ? reg_csr_3918 : _GEN_3917; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3919 = 12'hf4f == csr_addr[11:0] ? reg_csr_3919 : _GEN_3918; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3920 = 12'hf50 == csr_addr[11:0] ? reg_csr_3920 : _GEN_3919; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3921 = 12'hf51 == csr_addr[11:0] ? reg_csr_3921 : _GEN_3920; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3922 = 12'hf52 == csr_addr[11:0] ? reg_csr_3922 : _GEN_3921; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3923 = 12'hf53 == csr_addr[11:0] ? reg_csr_3923 : _GEN_3922; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3924 = 12'hf54 == csr_addr[11:0] ? reg_csr_3924 : _GEN_3923; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3925 = 12'hf55 == csr_addr[11:0] ? reg_csr_3925 : _GEN_3924; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3926 = 12'hf56 == csr_addr[11:0] ? reg_csr_3926 : _GEN_3925; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3927 = 12'hf57 == csr_addr[11:0] ? reg_csr_3927 : _GEN_3926; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3928 = 12'hf58 == csr_addr[11:0] ? reg_csr_3928 : _GEN_3927; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3929 = 12'hf59 == csr_addr[11:0] ? reg_csr_3929 : _GEN_3928; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3930 = 12'hf5a == csr_addr[11:0] ? reg_csr_3930 : _GEN_3929; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3931 = 12'hf5b == csr_addr[11:0] ? reg_csr_3931 : _GEN_3930; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3932 = 12'hf5c == csr_addr[11:0] ? reg_csr_3932 : _GEN_3931; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3933 = 12'hf5d == csr_addr[11:0] ? reg_csr_3933 : _GEN_3932; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3934 = 12'hf5e == csr_addr[11:0] ? reg_csr_3934 : _GEN_3933; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3935 = 12'hf5f == csr_addr[11:0] ? reg_csr_3935 : _GEN_3934; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3936 = 12'hf60 == csr_addr[11:0] ? reg_csr_3936 : _GEN_3935; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3937 = 12'hf61 == csr_addr[11:0] ? reg_csr_3937 : _GEN_3936; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3938 = 12'hf62 == csr_addr[11:0] ? reg_csr_3938 : _GEN_3937; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3939 = 12'hf63 == csr_addr[11:0] ? reg_csr_3939 : _GEN_3938; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3940 = 12'hf64 == csr_addr[11:0] ? reg_csr_3940 : _GEN_3939; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3941 = 12'hf65 == csr_addr[11:0] ? reg_csr_3941 : _GEN_3940; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3942 = 12'hf66 == csr_addr[11:0] ? reg_csr_3942 : _GEN_3941; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3943 = 12'hf67 == csr_addr[11:0] ? reg_csr_3943 : _GEN_3942; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3944 = 12'hf68 == csr_addr[11:0] ? reg_csr_3944 : _GEN_3943; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3945 = 12'hf69 == csr_addr[11:0] ? reg_csr_3945 : _GEN_3944; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3946 = 12'hf6a == csr_addr[11:0] ? reg_csr_3946 : _GEN_3945; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3947 = 12'hf6b == csr_addr[11:0] ? reg_csr_3947 : _GEN_3946; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3948 = 12'hf6c == csr_addr[11:0] ? reg_csr_3948 : _GEN_3947; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3949 = 12'hf6d == csr_addr[11:0] ? reg_csr_3949 : _GEN_3948; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3950 = 12'hf6e == csr_addr[11:0] ? reg_csr_3950 : _GEN_3949; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3951 = 12'hf6f == csr_addr[11:0] ? reg_csr_3951 : _GEN_3950; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3952 = 12'hf70 == csr_addr[11:0] ? reg_csr_3952 : _GEN_3951; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3953 = 12'hf71 == csr_addr[11:0] ? reg_csr_3953 : _GEN_3952; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3954 = 12'hf72 == csr_addr[11:0] ? reg_csr_3954 : _GEN_3953; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3955 = 12'hf73 == csr_addr[11:0] ? reg_csr_3955 : _GEN_3954; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3956 = 12'hf74 == csr_addr[11:0] ? reg_csr_3956 : _GEN_3955; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3957 = 12'hf75 == csr_addr[11:0] ? reg_csr_3957 : _GEN_3956; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3958 = 12'hf76 == csr_addr[11:0] ? reg_csr_3958 : _GEN_3957; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3959 = 12'hf77 == csr_addr[11:0] ? reg_csr_3959 : _GEN_3958; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3960 = 12'hf78 == csr_addr[11:0] ? reg_csr_3960 : _GEN_3959; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3961 = 12'hf79 == csr_addr[11:0] ? reg_csr_3961 : _GEN_3960; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3962 = 12'hf7a == csr_addr[11:0] ? reg_csr_3962 : _GEN_3961; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3963 = 12'hf7b == csr_addr[11:0] ? reg_csr_3963 : _GEN_3962; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3964 = 12'hf7c == csr_addr[11:0] ? reg_csr_3964 : _GEN_3963; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3965 = 12'hf7d == csr_addr[11:0] ? reg_csr_3965 : _GEN_3964; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3966 = 12'hf7e == csr_addr[11:0] ? reg_csr_3966 : _GEN_3965; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3967 = 12'hf7f == csr_addr[11:0] ? reg_csr_3967 : _GEN_3966; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3968 = 12'hf80 == csr_addr[11:0] ? reg_csr_3968 : _GEN_3967; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3969 = 12'hf81 == csr_addr[11:0] ? reg_csr_3969 : _GEN_3968; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3970 = 12'hf82 == csr_addr[11:0] ? reg_csr_3970 : _GEN_3969; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3971 = 12'hf83 == csr_addr[11:0] ? reg_csr_3971 : _GEN_3970; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3972 = 12'hf84 == csr_addr[11:0] ? reg_csr_3972 : _GEN_3971; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3973 = 12'hf85 == csr_addr[11:0] ? reg_csr_3973 : _GEN_3972; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3974 = 12'hf86 == csr_addr[11:0] ? reg_csr_3974 : _GEN_3973; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3975 = 12'hf87 == csr_addr[11:0] ? reg_csr_3975 : _GEN_3974; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3976 = 12'hf88 == csr_addr[11:0] ? reg_csr_3976 : _GEN_3975; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3977 = 12'hf89 == csr_addr[11:0] ? reg_csr_3977 : _GEN_3976; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3978 = 12'hf8a == csr_addr[11:0] ? reg_csr_3978 : _GEN_3977; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3979 = 12'hf8b == csr_addr[11:0] ? reg_csr_3979 : _GEN_3978; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3980 = 12'hf8c == csr_addr[11:0] ? reg_csr_3980 : _GEN_3979; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3981 = 12'hf8d == csr_addr[11:0] ? reg_csr_3981 : _GEN_3980; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3982 = 12'hf8e == csr_addr[11:0] ? reg_csr_3982 : _GEN_3981; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3983 = 12'hf8f == csr_addr[11:0] ? reg_csr_3983 : _GEN_3982; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3984 = 12'hf90 == csr_addr[11:0] ? reg_csr_3984 : _GEN_3983; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3985 = 12'hf91 == csr_addr[11:0] ? reg_csr_3985 : _GEN_3984; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3986 = 12'hf92 == csr_addr[11:0] ? reg_csr_3986 : _GEN_3985; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3987 = 12'hf93 == csr_addr[11:0] ? reg_csr_3987 : _GEN_3986; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3988 = 12'hf94 == csr_addr[11:0] ? reg_csr_3988 : _GEN_3987; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3989 = 12'hf95 == csr_addr[11:0] ? reg_csr_3989 : _GEN_3988; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3990 = 12'hf96 == csr_addr[11:0] ? reg_csr_3990 : _GEN_3989; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3991 = 12'hf97 == csr_addr[11:0] ? reg_csr_3991 : _GEN_3990; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3992 = 12'hf98 == csr_addr[11:0] ? reg_csr_3992 : _GEN_3991; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3993 = 12'hf99 == csr_addr[11:0] ? reg_csr_3993 : _GEN_3992; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3994 = 12'hf9a == csr_addr[11:0] ? reg_csr_3994 : _GEN_3993; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3995 = 12'hf9b == csr_addr[11:0] ? reg_csr_3995 : _GEN_3994; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3996 = 12'hf9c == csr_addr[11:0] ? reg_csr_3996 : _GEN_3995; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3997 = 12'hf9d == csr_addr[11:0] ? reg_csr_3997 : _GEN_3996; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3998 = 12'hf9e == csr_addr[11:0] ? reg_csr_3998 : _GEN_3997; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_3999 = 12'hf9f == csr_addr[11:0] ? reg_csr_3999 : _GEN_3998; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4000 = 12'hfa0 == csr_addr[11:0] ? reg_csr_4000 : _GEN_3999; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4001 = 12'hfa1 == csr_addr[11:0] ? reg_csr_4001 : _GEN_4000; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4002 = 12'hfa2 == csr_addr[11:0] ? reg_csr_4002 : _GEN_4001; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4003 = 12'hfa3 == csr_addr[11:0] ? reg_csr_4003 : _GEN_4002; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4004 = 12'hfa4 == csr_addr[11:0] ? reg_csr_4004 : _GEN_4003; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4005 = 12'hfa5 == csr_addr[11:0] ? reg_csr_4005 : _GEN_4004; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4006 = 12'hfa6 == csr_addr[11:0] ? reg_csr_4006 : _GEN_4005; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4007 = 12'hfa7 == csr_addr[11:0] ? reg_csr_4007 : _GEN_4006; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4008 = 12'hfa8 == csr_addr[11:0] ? reg_csr_4008 : _GEN_4007; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4009 = 12'hfa9 == csr_addr[11:0] ? reg_csr_4009 : _GEN_4008; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4010 = 12'hfaa == csr_addr[11:0] ? reg_csr_4010 : _GEN_4009; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4011 = 12'hfab == csr_addr[11:0] ? reg_csr_4011 : _GEN_4010; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4012 = 12'hfac == csr_addr[11:0] ? reg_csr_4012 : _GEN_4011; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4013 = 12'hfad == csr_addr[11:0] ? reg_csr_4013 : _GEN_4012; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4014 = 12'hfae == csr_addr[11:0] ? reg_csr_4014 : _GEN_4013; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4015 = 12'hfaf == csr_addr[11:0] ? reg_csr_4015 : _GEN_4014; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4016 = 12'hfb0 == csr_addr[11:0] ? reg_csr_4016 : _GEN_4015; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4017 = 12'hfb1 == csr_addr[11:0] ? reg_csr_4017 : _GEN_4016; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4018 = 12'hfb2 == csr_addr[11:0] ? reg_csr_4018 : _GEN_4017; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4019 = 12'hfb3 == csr_addr[11:0] ? reg_csr_4019 : _GEN_4018; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4020 = 12'hfb4 == csr_addr[11:0] ? reg_csr_4020 : _GEN_4019; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4021 = 12'hfb5 == csr_addr[11:0] ? reg_csr_4021 : _GEN_4020; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4022 = 12'hfb6 == csr_addr[11:0] ? reg_csr_4022 : _GEN_4021; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4023 = 12'hfb7 == csr_addr[11:0] ? reg_csr_4023 : _GEN_4022; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4024 = 12'hfb8 == csr_addr[11:0] ? reg_csr_4024 : _GEN_4023; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4025 = 12'hfb9 == csr_addr[11:0] ? reg_csr_4025 : _GEN_4024; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4026 = 12'hfba == csr_addr[11:0] ? reg_csr_4026 : _GEN_4025; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4027 = 12'hfbb == csr_addr[11:0] ? reg_csr_4027 : _GEN_4026; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4028 = 12'hfbc == csr_addr[11:0] ? reg_csr_4028 : _GEN_4027; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4029 = 12'hfbd == csr_addr[11:0] ? reg_csr_4029 : _GEN_4028; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4030 = 12'hfbe == csr_addr[11:0] ? reg_csr_4030 : _GEN_4029; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4031 = 12'hfbf == csr_addr[11:0] ? reg_csr_4031 : _GEN_4030; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4032 = 12'hfc0 == csr_addr[11:0] ? reg_csr_4032 : _GEN_4031; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4033 = 12'hfc1 == csr_addr[11:0] ? reg_csr_4033 : _GEN_4032; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4034 = 12'hfc2 == csr_addr[11:0] ? reg_csr_4034 : _GEN_4033; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4035 = 12'hfc3 == csr_addr[11:0] ? reg_csr_4035 : _GEN_4034; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4036 = 12'hfc4 == csr_addr[11:0] ? reg_csr_4036 : _GEN_4035; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4037 = 12'hfc5 == csr_addr[11:0] ? reg_csr_4037 : _GEN_4036; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4038 = 12'hfc6 == csr_addr[11:0] ? reg_csr_4038 : _GEN_4037; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4039 = 12'hfc7 == csr_addr[11:0] ? reg_csr_4039 : _GEN_4038; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4040 = 12'hfc8 == csr_addr[11:0] ? reg_csr_4040 : _GEN_4039; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4041 = 12'hfc9 == csr_addr[11:0] ? reg_csr_4041 : _GEN_4040; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4042 = 12'hfca == csr_addr[11:0] ? reg_csr_4042 : _GEN_4041; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4043 = 12'hfcb == csr_addr[11:0] ? reg_csr_4043 : _GEN_4042; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4044 = 12'hfcc == csr_addr[11:0] ? reg_csr_4044 : _GEN_4043; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4045 = 12'hfcd == csr_addr[11:0] ? reg_csr_4045 : _GEN_4044; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4046 = 12'hfce == csr_addr[11:0] ? reg_csr_4046 : _GEN_4045; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4047 = 12'hfcf == csr_addr[11:0] ? reg_csr_4047 : _GEN_4046; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4048 = 12'hfd0 == csr_addr[11:0] ? reg_csr_4048 : _GEN_4047; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4049 = 12'hfd1 == csr_addr[11:0] ? reg_csr_4049 : _GEN_4048; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4050 = 12'hfd2 == csr_addr[11:0] ? reg_csr_4050 : _GEN_4049; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4051 = 12'hfd3 == csr_addr[11:0] ? reg_csr_4051 : _GEN_4050; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4052 = 12'hfd4 == csr_addr[11:0] ? reg_csr_4052 : _GEN_4051; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4053 = 12'hfd5 == csr_addr[11:0] ? reg_csr_4053 : _GEN_4052; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4054 = 12'hfd6 == csr_addr[11:0] ? reg_csr_4054 : _GEN_4053; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4055 = 12'hfd7 == csr_addr[11:0] ? reg_csr_4055 : _GEN_4054; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4056 = 12'hfd8 == csr_addr[11:0] ? reg_csr_4056 : _GEN_4055; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4057 = 12'hfd9 == csr_addr[11:0] ? reg_csr_4057 : _GEN_4056; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4058 = 12'hfda == csr_addr[11:0] ? reg_csr_4058 : _GEN_4057; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4059 = 12'hfdb == csr_addr[11:0] ? reg_csr_4059 : _GEN_4058; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4060 = 12'hfdc == csr_addr[11:0] ? reg_csr_4060 : _GEN_4059; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4061 = 12'hfdd == csr_addr[11:0] ? reg_csr_4061 : _GEN_4060; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4062 = 12'hfde == csr_addr[11:0] ? reg_csr_4062 : _GEN_4061; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4063 = 12'hfdf == csr_addr[11:0] ? reg_csr_4063 : _GEN_4062; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4064 = 12'hfe0 == csr_addr[11:0] ? reg_csr_4064 : _GEN_4063; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4065 = 12'hfe1 == csr_addr[11:0] ? reg_csr_4065 : _GEN_4064; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4066 = 12'hfe2 == csr_addr[11:0] ? reg_csr_4066 : _GEN_4065; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4067 = 12'hfe3 == csr_addr[11:0] ? reg_csr_4067 : _GEN_4066; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4068 = 12'hfe4 == csr_addr[11:0] ? reg_csr_4068 : _GEN_4067; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4069 = 12'hfe5 == csr_addr[11:0] ? reg_csr_4069 : _GEN_4068; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4070 = 12'hfe6 == csr_addr[11:0] ? reg_csr_4070 : _GEN_4069; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4071 = 12'hfe7 == csr_addr[11:0] ? reg_csr_4071 : _GEN_4070; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4072 = 12'hfe8 == csr_addr[11:0] ? reg_csr_4072 : _GEN_4071; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4073 = 12'hfe9 == csr_addr[11:0] ? reg_csr_4073 : _GEN_4072; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4074 = 12'hfea == csr_addr[11:0] ? reg_csr_4074 : _GEN_4073; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4075 = 12'hfeb == csr_addr[11:0] ? reg_csr_4075 : _GEN_4074; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4076 = 12'hfec == csr_addr[11:0] ? reg_csr_4076 : _GEN_4075; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4077 = 12'hfed == csr_addr[11:0] ? reg_csr_4077 : _GEN_4076; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4078 = 12'hfee == csr_addr[11:0] ? reg_csr_4078 : _GEN_4077; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4079 = 12'hfef == csr_addr[11:0] ? reg_csr_4079 : _GEN_4078; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4080 = 12'hff0 == csr_addr[11:0] ? reg_csr_4080 : _GEN_4079; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4081 = 12'hff1 == csr_addr[11:0] ? reg_csr_4081 : _GEN_4080; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4082 = 12'hff2 == csr_addr[11:0] ? reg_csr_4082 : _GEN_4081; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4083 = 12'hff3 == csr_addr[11:0] ? reg_csr_4083 : _GEN_4082; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4084 = 12'hff4 == csr_addr[11:0] ? reg_csr_4084 : _GEN_4083; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4085 = 12'hff5 == csr_addr[11:0] ? reg_csr_4085 : _GEN_4084; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4086 = 12'hff6 == csr_addr[11:0] ? reg_csr_4086 : _GEN_4085; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4087 = 12'hff7 == csr_addr[11:0] ? reg_csr_4087 : _GEN_4086; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4088 = 12'hff8 == csr_addr[11:0] ? reg_csr_4088 : _GEN_4087; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4089 = 12'hff9 == csr_addr[11:0] ? reg_csr_4089 : _GEN_4088; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4090 = 12'hffa == csr_addr[11:0] ? reg_csr_4090 : _GEN_4089; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4091 = 12'hffb == csr_addr[11:0] ? reg_csr_4091 : _GEN_4090; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4092 = 12'hffc == csr_addr[11:0] ? reg_csr_4092 : _GEN_4091; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4093 = 12'hffd == csr_addr[11:0] ? reg_csr_4093 : _GEN_4092; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4094 = 12'hffe == csr_addr[11:0] ? reg_csr_4094 : _GEN_4093; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _GEN_4095 = 12'hfff == csr_addr[11:0] ? reg_csr_4095 : _GEN_4094; // @[CSR.scala 45:43 CSR.scala 45:43]
  wire [31:0] _csr_wdata_T_2 = _GEN_4095 | io_in_id_io_op1_data; // @[CSR.scala 45:43]
  wire  _csr_wdata_T_3 = io_in_id_io_csr_cmd == 3'h3; // @[CSR.scala 46:18]
  wire [31:0] _csr_wdata_T_4 = ~io_in_id_io_op1_data; // @[CSR.scala 46:45]
  wire [31:0] _csr_wdata_T_5 = _GEN_4095 & _csr_wdata_T_4; // @[CSR.scala 46:43]
  wire [31:0] _csr_wdata_T_7 = _csr_addr_T ? 32'hb : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _csr_wdata_T_8 = _csr_wdata_T_3 ? _csr_wdata_T_5 : _csr_wdata_T_7; // @[Mux.scala 98:16]
  wire [31:0] _csr_wdata_T_9 = _csr_wdata_T_1 ? _csr_wdata_T_2 : _csr_wdata_T_8; // @[Mux.scala 98:16]
  wire [31:0] csr_wdata = _csr_wdata_T ? io_in_id_io_op1_data : _csr_wdata_T_9; // @[Mux.scala 98:16]
  wire  _T_3 = ~reset; // @[CSR.scala 58:11]
  assign io_out_csr_rdata = 12'hfff == csr_addr[11:0] ? reg_csr_4095 : _GEN_4094; // @[CSR.scala 45:43 CSR.scala 45:43]
  assign io_out_trap_vector = reg_csr_773; // @[CSR.scala 55:25]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_0 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_0 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_0 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_5 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_5 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_5 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_6 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_6 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_6 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_7 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_7 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_7 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_8 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_8 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_8 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_9 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_9 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_9 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_10 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_10 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_10 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_11 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_11 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_11 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_12 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_12 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_12 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_13 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_13 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_13 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_14 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_14 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_14 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_15 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_15 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_15 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_16 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_16 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_16 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_17 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_17 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_17 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_18 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_18 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_18 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_19 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_19 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_19 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_20 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_20 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_20 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_21 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_21 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_21 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_22 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_22 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_22 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_23 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_23 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_23 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_24 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_24 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_24 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_25 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_25 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_25 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_26 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_26 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_26 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_27 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_27 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_27 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_28 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_28 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_28 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_29 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_29 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_29 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_30 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_30 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_30 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_31 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_31 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_31 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_32 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_32 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_32 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_33 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_33 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_33 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_34 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_34 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_34 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_35 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_35 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_35 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_36 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_36 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_36 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_37 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_37 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_37 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_38 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_38 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_38 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_39 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_39 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_39 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_40 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_40 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_40 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_41 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_41 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_41 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_42 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_42 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_42 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_43 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_43 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_43 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_44 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_44 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_44 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_45 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_45 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_45 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_46 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_46 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_46 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_47 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_47 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_47 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_48 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_48 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_48 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_49 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_49 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_49 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_50 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_50 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_50 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_51 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_51 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_51 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_52 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_52 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_52 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_53 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_53 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_53 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_54 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_54 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_54 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_55 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_55 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_55 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_56 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_56 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_56 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_57 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_57 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_57 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_58 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_58 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_58 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_59 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_59 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_59 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_60 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_60 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_60 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_61 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_61 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_61 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_62 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_62 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_62 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_63 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_63 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_63 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_64 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_64 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_64 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_65 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_65 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_65 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_66 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_66 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_66 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_67 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_67 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_67 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_68 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_68 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_68 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_69 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_69 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_69 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_70 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_70 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_70 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_71 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_71 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_71 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_72 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_72 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_72 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_73 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_73 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_73 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_74 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_74 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_74 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_75 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_75 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_75 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_76 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_76 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_76 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_77 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_77 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_77 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_78 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_78 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_78 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_79 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_79 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_79 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_80 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_80 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_80 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_81 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_81 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_81 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_82 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_82 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_82 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_83 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_83 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_83 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_84 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_84 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_84 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_85 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_85 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_85 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_86 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_86 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_86 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_87 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_87 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_87 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_88 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_88 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_88 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_89 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_89 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_89 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_90 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_90 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_90 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_91 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_91 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_91 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_92 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_92 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_92 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_93 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_93 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_93 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_94 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_94 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_94 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_95 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_95 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_95 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_96 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_96 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_96 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_97 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_97 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_97 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_98 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_98 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_98 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_99 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_99 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_99 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_100 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_100 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_100 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_101 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_101 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_101 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_102 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_102 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_102 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_103 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_103 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_103 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_104 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_104 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_104 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_105 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_105 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_105 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_106 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_106 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_106 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_107 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_107 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_107 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_108 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_108 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_108 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_109 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_109 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_109 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_110 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_110 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_110 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_111 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_111 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_111 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_112 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_112 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_112 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_113 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_113 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_113 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_114 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_114 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_114 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_115 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_115 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_115 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_116 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_116 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_116 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_117 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_117 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_117 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_118 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_118 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_118 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_119 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_119 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_119 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_120 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_120 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_120 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_121 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_121 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_121 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_122 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_122 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_122 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_123 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_123 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_123 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_124 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_124 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_124 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_125 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_125 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_125 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_126 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_126 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_126 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_127 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_127 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_127 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_128 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_128 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_128 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_129 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_129 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_129 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_130 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_130 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_130 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_131 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_131 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_131 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_132 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_132 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_132 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_133 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_133 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_133 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_134 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_134 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_134 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_135 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_135 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_135 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_136 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_136 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_136 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_137 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_137 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_137 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_138 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_138 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_138 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_139 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_139 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_139 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_140 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_140 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_140 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_141 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_141 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_141 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_142 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_142 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_142 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_143 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_143 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_143 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_144 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_144 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_144 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_145 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_145 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_145 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_146 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_146 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_146 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_147 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_147 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_147 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_148 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_148 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_148 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_149 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_149 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_149 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_150 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_150 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_150 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_151 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_151 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_151 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_152 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_152 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_152 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_153 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_153 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_153 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_154 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_154 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_154 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_155 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_155 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_155 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_156 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_156 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_156 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_157 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_157 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_157 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_158 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_158 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_158 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_159 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_159 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_159 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_160 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_160 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_160 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_161 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_161 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_161 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_162 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_162 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_162 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_163 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_163 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_163 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_164 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_164 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_164 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_165 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_165 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_165 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_166 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_166 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_166 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_167 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_167 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_167 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_168 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_168 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_168 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_169 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_169 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_169 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_170 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_170 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_170 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_171 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_171 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_171 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_172 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_172 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_172 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_173 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_173 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_173 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_174 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_174 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_174 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_175 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_175 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_175 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_176 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_176 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_176 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_177 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_177 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_177 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_178 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_178 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_178 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_179 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_179 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_179 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_180 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_180 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_180 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_181 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_181 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_181 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_182 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_182 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_182 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_183 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_183 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_183 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_184 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_184 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_184 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_185 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_185 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_185 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_186 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_186 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_186 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_187 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_187 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_187 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_188 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_188 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_188 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_189 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_189 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_189 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_190 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_190 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_190 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_191 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_191 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_191 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_192 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_192 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_192 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_193 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_193 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_193 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_194 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_194 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_194 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_195 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_195 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_195 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_196 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_196 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_196 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_197 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_197 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_197 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_198 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_198 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_198 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_199 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_199 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_199 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_200 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_200 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_200 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_201 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_201 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_201 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_202 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_202 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_202 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_203 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_203 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_203 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_204 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_204 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_204 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_205 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_205 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_205 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_206 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_206 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_206 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_207 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_207 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_207 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_208 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_208 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_208 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_209 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_209 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_209 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_210 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_210 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_210 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_211 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_211 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_211 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_212 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_212 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_212 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_213 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_213 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_213 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_214 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_214 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_214 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_215 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_215 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_215 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_216 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_216 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_216 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_217 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_217 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_217 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_218 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_218 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_218 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_219 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_219 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_219 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_220 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_220 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_220 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_221 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_221 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_221 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_222 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_222 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_222 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_223 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_223 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_223 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_224 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_224 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_224 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_225 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_225 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_225 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_226 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_226 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_226 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_227 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_227 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_227 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_228 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_228 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_228 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_229 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_229 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_229 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_230 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_230 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_230 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_231 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_231 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_231 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_232 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_232 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_232 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_233 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_233 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_233 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_234 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_234 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_234 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_235 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_235 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_235 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_236 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_236 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_236 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_237 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_237 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_237 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_238 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_238 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_238 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_239 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_239 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_239 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_240 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_240 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_240 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_241 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_241 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_241 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_242 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_242 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_242 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_243 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_243 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_243 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_244 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_244 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_244 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_245 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_245 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_245 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_246 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_246 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_246 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_247 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_247 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_247 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_248 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_248 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_248 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_249 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_249 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_249 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_250 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_250 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_250 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_251 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_251 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_251 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_252 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_252 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_252 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_253 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_253 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_253 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_254 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_254 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_254 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_255 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_255 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_255 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_256 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h100 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_256 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_256 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_257 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h101 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_257 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_257 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_258 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h102 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_258 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_258 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_259 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h103 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_259 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_259 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_260 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h104 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_260 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_260 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_261 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h105 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_261 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_261 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_262 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h106 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_262 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_262 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_263 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h107 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_263 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_263 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_264 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h108 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_264 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_264 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_265 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h109 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_265 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_265 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_266 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_266 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_266 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_267 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_267 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_267 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_268 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_268 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_268 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_269 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_269 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_269 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_270 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_270 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_270 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_271 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h10f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_271 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_271 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_272 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h110 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_272 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_272 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_273 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h111 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_273 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_273 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_274 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h112 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_274 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_274 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_275 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h113 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_275 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_275 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_276 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h114 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_276 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_276 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_277 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h115 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_277 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_277 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_278 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h116 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_278 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_278 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_279 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h117 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_279 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_279 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_280 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h118 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_280 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_280 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_281 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h119 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_281 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_281 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_282 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_282 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_282 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_283 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_283 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_283 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_284 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_284 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_284 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_285 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_285 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_285 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_286 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_286 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_286 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_287 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h11f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_287 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_287 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_288 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h120 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_288 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_288 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_289 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h121 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_289 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_289 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_290 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h122 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_290 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_290 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_291 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h123 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_291 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_291 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_292 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h124 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_292 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_292 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_293 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h125 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_293 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_293 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_294 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h126 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_294 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_294 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_295 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h127 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_295 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_295 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_296 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h128 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_296 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_296 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_297 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h129 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_297 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_297 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_298 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_298 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_298 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_299 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_299 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_299 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_300 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_300 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_300 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_301 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_301 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_301 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_302 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_302 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_302 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_303 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h12f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_303 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_303 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_304 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h130 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_304 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_304 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_305 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h131 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_305 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_305 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_306 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h132 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_306 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_306 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_307 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h133 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_307 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_307 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_308 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h134 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_308 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_308 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_309 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h135 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_309 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_309 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_310 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h136 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_310 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_310 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_311 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h137 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_311 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_311 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_312 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h138 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_312 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_312 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_313 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h139 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_313 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_313 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_314 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_314 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_314 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_315 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_315 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_315 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_316 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_316 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_316 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_317 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_317 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_317 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_318 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_318 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_318 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_319 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h13f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_319 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_319 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_320 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h140 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_320 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_320 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_321 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h141 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_321 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_321 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_322 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h142 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_322 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_322 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_323 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h143 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_323 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_323 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_324 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h144 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_324 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_324 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_325 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h145 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_325 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_325 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_326 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h146 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_326 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_326 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_327 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h147 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_327 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_327 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_328 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h148 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_328 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_328 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_329 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h149 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_329 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_329 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_330 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_330 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_330 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_331 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_331 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_331 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_332 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_332 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_332 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_333 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_333 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_333 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_334 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_334 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_334 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_335 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h14f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_335 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_335 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_336 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h150 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_336 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_336 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_337 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h151 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_337 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_337 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_338 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h152 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_338 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_338 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_339 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h153 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_339 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_339 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_340 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h154 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_340 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_340 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_341 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h155 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_341 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_341 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_342 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h156 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_342 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_342 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_343 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h157 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_343 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_343 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_344 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h158 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_344 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_344 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_345 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h159 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_345 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_345 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_346 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_346 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_346 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_347 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_347 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_347 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_348 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_348 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_348 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_349 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_349 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_349 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_350 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_350 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_350 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_351 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h15f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_351 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_351 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_352 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h160 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_352 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_352 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_353 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h161 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_353 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_353 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_354 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h162 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_354 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_354 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_355 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h163 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_355 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_355 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_356 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h164 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_356 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_356 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_357 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h165 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_357 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_357 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_358 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h166 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_358 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_358 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_359 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h167 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_359 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_359 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_360 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h168 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_360 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_360 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_361 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h169 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_361 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_361 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_362 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_362 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_362 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_363 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_363 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_363 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_364 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_364 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_364 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_365 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_365 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_365 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_366 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_366 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_366 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_367 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h16f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_367 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_367 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_368 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h170 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_368 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_368 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_369 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h171 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_369 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_369 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_370 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h172 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_370 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_370 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_371 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h173 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_371 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_371 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_372 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h174 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_372 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_372 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_373 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h175 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_373 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_373 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_374 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h176 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_374 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_374 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_375 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h177 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_375 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_375 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_376 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h178 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_376 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_376 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_377 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h179 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_377 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_377 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_378 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_378 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_378 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_379 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_379 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_379 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_380 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_380 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_380 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_381 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_381 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_381 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_382 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_382 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_382 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_383 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h17f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_383 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_383 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_384 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h180 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_384 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_384 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_385 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h181 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_385 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_385 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_386 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h182 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_386 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_386 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_387 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h183 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_387 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_387 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_388 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h184 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_388 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_388 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_389 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h185 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_389 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_389 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_390 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h186 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_390 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_390 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_391 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h187 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_391 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_391 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_392 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h188 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_392 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_392 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_393 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h189 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_393 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_393 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_394 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_394 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_394 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_395 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_395 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_395 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_396 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_396 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_396 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_397 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_397 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_397 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_398 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_398 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_398 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_399 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h18f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_399 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_399 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_400 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h190 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_400 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_400 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_401 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h191 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_401 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_401 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_402 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h192 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_402 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_402 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_403 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h193 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_403 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_403 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_404 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h194 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_404 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_404 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_405 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h195 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_405 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_405 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_406 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h196 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_406 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_406 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_407 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h197 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_407 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_407 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_408 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h198 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_408 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_408 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_409 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h199 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_409 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_409 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_410 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_410 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_410 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_411 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_411 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_411 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_412 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_412 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_412 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_413 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_413 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_413 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_414 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_414 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_414 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_415 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h19f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_415 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_415 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_416 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_416 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_416 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_417 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_417 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_417 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_418 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_418 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_418 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_419 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_419 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_419 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_420 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_420 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_420 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_421 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_421 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_421 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_422 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_422 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_422 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_423 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_423 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_423 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_424 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_424 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_424 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_425 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_425 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_425 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_426 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_426 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_426 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_427 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_427 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_427 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_428 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_428 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_428 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_429 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_429 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_429 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_430 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_430 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_430 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_431 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_431 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_431 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_432 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_432 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_432 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_433 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_433 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_433 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_434 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_434 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_434 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_435 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_435 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_435 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_436 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_436 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_436 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_437 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_437 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_437 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_438 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_438 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_438 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_439 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_439 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_439 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_440 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_440 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_440 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_441 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_441 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_441 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_442 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_442 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_442 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_443 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_443 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_443 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_444 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_444 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_444 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_445 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_445 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_445 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_446 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_446 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_446 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_447 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_447 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_447 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_448 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_448 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_448 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_449 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_449 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_449 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_450 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_450 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_450 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_451 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_451 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_451 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_452 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_452 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_452 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_453 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_453 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_453 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_454 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_454 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_454 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_455 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_455 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_455 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_456 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_456 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_456 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_457 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_457 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_457 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_458 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_458 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_458 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_459 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_459 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_459 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_460 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_460 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_460 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_461 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_461 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_461 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_462 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_462 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_462 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_463 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_463 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_463 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_464 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_464 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_464 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_465 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_465 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_465 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_466 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_466 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_466 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_467 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_467 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_467 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_468 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_468 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_468 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_469 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_469 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_469 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_470 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_470 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_470 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_471 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_471 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_471 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_472 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_472 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_472 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_473 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_473 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_473 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_474 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_474 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_474 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_475 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_475 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_475 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_476 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_476 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_476 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_477 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_477 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_477 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_478 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_478 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_478 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_479 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_479 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_479 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_480 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_480 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_480 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_481 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_481 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_481 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_482 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_482 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_482 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_483 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_483 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_483 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_484 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_484 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_484 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_485 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_485 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_485 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_486 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_486 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_486 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_487 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_487 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_487 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_488 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_488 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_488 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_489 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_489 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_489 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_490 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_490 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_490 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_491 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_491 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_491 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_492 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_492 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_492 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_493 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_493 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_493 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_494 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_494 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_494 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_495 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_495 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_495 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_496 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_496 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_496 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_497 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_497 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_497 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_498 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_498 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_498 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_499 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_499 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_499 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_500 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_500 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_500 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_501 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_501 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_501 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_502 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_502 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_502 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_503 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_503 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_503 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_504 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_504 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_504 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_505 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_505 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_505 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_506 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_506 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_506 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_507 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_507 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_507 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_508 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_508 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_508 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_509 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_509 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_509 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_510 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_510 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_510 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_511 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h1ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_511 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_511 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_512 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h200 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_512 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_512 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_513 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h201 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_513 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_513 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_514 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h202 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_514 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_514 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_515 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h203 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_515 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_515 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_516 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h204 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_516 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_516 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_517 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h205 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_517 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_517 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_518 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h206 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_518 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_518 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_519 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h207 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_519 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_519 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_520 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h208 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_520 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_520 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_521 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h209 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_521 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_521 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_522 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_522 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_522 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_523 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_523 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_523 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_524 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_524 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_524 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_525 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_525 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_525 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_526 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_526 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_526 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_527 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h20f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_527 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_527 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_528 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h210 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_528 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_528 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_529 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h211 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_529 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_529 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_530 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h212 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_530 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_530 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_531 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h213 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_531 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_531 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_532 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h214 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_532 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_532 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_533 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h215 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_533 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_533 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_534 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h216 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_534 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_534 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_535 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h217 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_535 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_535 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_536 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h218 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_536 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_536 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_537 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h219 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_537 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_537 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_538 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_538 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_538 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_539 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_539 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_539 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_540 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_540 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_540 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_541 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_541 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_541 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_542 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_542 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_542 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_543 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h21f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_543 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_543 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_544 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h220 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_544 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_544 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_545 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h221 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_545 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_545 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_546 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h222 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_546 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_546 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_547 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h223 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_547 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_547 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_548 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h224 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_548 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_548 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_549 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h225 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_549 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_549 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_550 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h226 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_550 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_550 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_551 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h227 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_551 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_551 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_552 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h228 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_552 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_552 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_553 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h229 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_553 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_553 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_554 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_554 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_554 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_555 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_555 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_555 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_556 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_556 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_556 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_557 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_557 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_557 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_558 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_558 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_558 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_559 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h22f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_559 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_559 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_560 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h230 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_560 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_560 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_561 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h231 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_561 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_561 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_562 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h232 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_562 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_562 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_563 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h233 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_563 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_563 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_564 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h234 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_564 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_564 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_565 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h235 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_565 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_565 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_566 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h236 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_566 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_566 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_567 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h237 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_567 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_567 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_568 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h238 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_568 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_568 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_569 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h239 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_569 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_569 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_570 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_570 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_570 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_571 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_571 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_571 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_572 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_572 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_572 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_573 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_573 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_573 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_574 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_574 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_574 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_575 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h23f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_575 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_575 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_576 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h240 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_576 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_576 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_577 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h241 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_577 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_577 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_578 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h242 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_578 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_578 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_579 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h243 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_579 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_579 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_580 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h244 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_580 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_580 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_581 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h245 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_581 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_581 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_582 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h246 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_582 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_582 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_583 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h247 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_583 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_583 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_584 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h248 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_584 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_584 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_585 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h249 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_585 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_585 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_586 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_586 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_586 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_587 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_587 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_587 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_588 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_588 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_588 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_589 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_589 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_589 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_590 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_590 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_590 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_591 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h24f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_591 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_591 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_592 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h250 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_592 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_592 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_593 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h251 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_593 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_593 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_594 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h252 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_594 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_594 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_595 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h253 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_595 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_595 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_596 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h254 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_596 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_596 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_597 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h255 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_597 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_597 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_598 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h256 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_598 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_598 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_599 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h257 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_599 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_599 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_600 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h258 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_600 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_600 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_601 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h259 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_601 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_601 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_602 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_602 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_602 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_603 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_603 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_603 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_604 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_604 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_604 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_605 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_605 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_605 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_606 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_606 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_606 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_607 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h25f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_607 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_607 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_608 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h260 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_608 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_608 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_609 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h261 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_609 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_609 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_610 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h262 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_610 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_610 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_611 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h263 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_611 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_611 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_612 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h264 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_612 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_612 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_613 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h265 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_613 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_613 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_614 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h266 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_614 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_614 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_615 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h267 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_615 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_615 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_616 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h268 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_616 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_616 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_617 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h269 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_617 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_617 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_618 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_618 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_618 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_619 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_619 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_619 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_620 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_620 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_620 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_621 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_621 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_621 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_622 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_622 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_622 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_623 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h26f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_623 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_623 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_624 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h270 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_624 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_624 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_625 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h271 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_625 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_625 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_626 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h272 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_626 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_626 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_627 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h273 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_627 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_627 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_628 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h274 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_628 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_628 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_629 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h275 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_629 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_629 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_630 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h276 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_630 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_630 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_631 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h277 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_631 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_631 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_632 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h278 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_632 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_632 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_633 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h279 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_633 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_633 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_634 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_634 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_634 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_635 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_635 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_635 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_636 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_636 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_636 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_637 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_637 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_637 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_638 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_638 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_638 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_639 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h27f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_639 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_639 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_640 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h280 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_640 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_640 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_641 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h281 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_641 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_641 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_642 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h282 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_642 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_642 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_643 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h283 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_643 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_643 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_644 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h284 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_644 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_644 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_645 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h285 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_645 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_645 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_646 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h286 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_646 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_646 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_647 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h287 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_647 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_647 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_648 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h288 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_648 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_648 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_649 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h289 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_649 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_649 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_650 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_650 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_650 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_651 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_651 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_651 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_652 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_652 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_652 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_653 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_653 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_653 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_654 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_654 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_654 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_655 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h28f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_655 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_655 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_656 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h290 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_656 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_656 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_657 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h291 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_657 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_657 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_658 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h292 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_658 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_658 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_659 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h293 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_659 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_659 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_660 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h294 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_660 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_660 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_661 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h295 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_661 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_661 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_662 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h296 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_662 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_662 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_663 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h297 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_663 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_663 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_664 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h298 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_664 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_664 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_665 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h299 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_665 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_665 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_666 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_666 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_666 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_667 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_667 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_667 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_668 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_668 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_668 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_669 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_669 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_669 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_670 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_670 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_670 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_671 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h29f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_671 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_671 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_672 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_672 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_672 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_673 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_673 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_673 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_674 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_674 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_674 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_675 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_675 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_675 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_676 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_676 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_676 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_677 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_677 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_677 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_678 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_678 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_678 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_679 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_679 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_679 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_680 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_680 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_680 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_681 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_681 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_681 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_682 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_682 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_682 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_683 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_683 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_683 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_684 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_684 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_684 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_685 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_685 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_685 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_686 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_686 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_686 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_687 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_687 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_687 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_688 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_688 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_688 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_689 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_689 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_689 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_690 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_690 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_690 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_691 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_691 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_691 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_692 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_692 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_692 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_693 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_693 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_693 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_694 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_694 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_694 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_695 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_695 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_695 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_696 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_696 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_696 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_697 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_697 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_697 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_698 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_698 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_698 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_699 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_699 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_699 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_700 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_700 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_700 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_701 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_701 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_701 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_702 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_702 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_702 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_703 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_703 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_703 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_704 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_704 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_704 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_705 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_705 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_705 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_706 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_706 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_706 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_707 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_707 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_707 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_708 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_708 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_708 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_709 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_709 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_709 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_710 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_710 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_710 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_711 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_711 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_711 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_712 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_712 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_712 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_713 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_713 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_713 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_714 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_714 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_714 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_715 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_715 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_715 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_716 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_716 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_716 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_717 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_717 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_717 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_718 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_718 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_718 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_719 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_719 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_719 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_720 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_720 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_720 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_721 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_721 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_721 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_722 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_722 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_722 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_723 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_723 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_723 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_724 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_724 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_724 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_725 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_725 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_725 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_726 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_726 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_726 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_727 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_727 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_727 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_728 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_728 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_728 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_729 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_729 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_729 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_730 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_730 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_730 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_731 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_731 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_731 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_732 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_732 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_732 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_733 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_733 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_733 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_734 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_734 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_734 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_735 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_735 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_735 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_736 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_736 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_736 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_737 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_737 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_737 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_738 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_738 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_738 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_739 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_739 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_739 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_740 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_740 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_740 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_741 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_741 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_741 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_742 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_742 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_742 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_743 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_743 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_743 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_744 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_744 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_744 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_745 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_745 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_745 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_746 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_746 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_746 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_747 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_747 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_747 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_748 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_748 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_748 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_749 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_749 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_749 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_750 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_750 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_750 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_751 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_751 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_751 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_752 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_752 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_752 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_753 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_753 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_753 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_754 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_754 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_754 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_755 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_755 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_755 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_756 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_756 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_756 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_757 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_757 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_757 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_758 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_758 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_758 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_759 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_759 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_759 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_760 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_760 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_760 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_761 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_761 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_761 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_762 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_762 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_762 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_763 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_763 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_763 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_764 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_764 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_764 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_765 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_765 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_765 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_766 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_766 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_766 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_767 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h2ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_767 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_767 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_768 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h300 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_768 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_768 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_769 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h301 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_769 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_769 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_770 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h302 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_770 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_770 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_771 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h303 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_771 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_771 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_772 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h304 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_772 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_772 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_773 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h305 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_773 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_773 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_774 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h306 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_774 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_774 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_775 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h307 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_775 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_775 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_776 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h308 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_776 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_776 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_777 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h309 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_777 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_777 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_778 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_778 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_778 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_779 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_779 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_779 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_780 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_780 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_780 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_781 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_781 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_781 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_782 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_782 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_782 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_783 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h30f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_783 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_783 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_784 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h310 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_784 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_784 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_785 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h311 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_785 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_785 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_786 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h312 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_786 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_786 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_787 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h313 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_787 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_787 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_788 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h314 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_788 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_788 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_789 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h315 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_789 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_789 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_790 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h316 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_790 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_790 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_791 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h317 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_791 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_791 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_792 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h318 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_792 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_792 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_793 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h319 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_793 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_793 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_794 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_794 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_794 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_795 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_795 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_795 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_796 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_796 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_796 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_797 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_797 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_797 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_798 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_798 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_798 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_799 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h31f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_799 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_799 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_800 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h320 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_800 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_800 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_801 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h321 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_801 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_801 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_802 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h322 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_802 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_802 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_803 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h323 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_803 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_803 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_804 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h324 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_804 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_804 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_805 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h325 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_805 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_805 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_806 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h326 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_806 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_806 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_807 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h327 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_807 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_807 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_808 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h328 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_808 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_808 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_809 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h329 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_809 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_809 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_810 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_810 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_810 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_811 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_811 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_811 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_812 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_812 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_812 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_813 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_813 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_813 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_814 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_814 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_814 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_815 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h32f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_815 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_815 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_816 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h330 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_816 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_816 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_817 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h331 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_817 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_817 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_818 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h332 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_818 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_818 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_819 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h333 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_819 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_819 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_820 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h334 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_820 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_820 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_821 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h335 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_821 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_821 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_822 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h336 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_822 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_822 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_823 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h337 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_823 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_823 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_824 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h338 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_824 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_824 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_825 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h339 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_825 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_825 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_826 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_826 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_826 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_827 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_827 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_827 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_828 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_828 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_828 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_829 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_829 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_829 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_830 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_830 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_830 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_831 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h33f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_831 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_831 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_832 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h340 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_832 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_832 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_833 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h341 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_833 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_833 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_834 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h342 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_834 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_834 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_835 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h343 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_835 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_835 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_836 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h344 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_836 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_836 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_837 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h345 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_837 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_837 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_838 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h346 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_838 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_838 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_839 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h347 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_839 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_839 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_840 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h348 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_840 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_840 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_841 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h349 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_841 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_841 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_842 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_842 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_842 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_843 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_843 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_843 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_844 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_844 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_844 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_845 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_845 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_845 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_846 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_846 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_846 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_847 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h34f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_847 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_847 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_848 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h350 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_848 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_848 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_849 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h351 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_849 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_849 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_850 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h352 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_850 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_850 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_851 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h353 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_851 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_851 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_852 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h354 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_852 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_852 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_853 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h355 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_853 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_853 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_854 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h356 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_854 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_854 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_855 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h357 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_855 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_855 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_856 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h358 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_856 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_856 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_857 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h359 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_857 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_857 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_858 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_858 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_858 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_859 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_859 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_859 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_860 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_860 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_860 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_861 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_861 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_861 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_862 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_862 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_862 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_863 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h35f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_863 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_863 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_864 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h360 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_864 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_864 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_865 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h361 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_865 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_865 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_866 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h362 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_866 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_866 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_867 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h363 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_867 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_867 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_868 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h364 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_868 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_868 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_869 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h365 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_869 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_869 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_870 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h366 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_870 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_870 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_871 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h367 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_871 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_871 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_872 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h368 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_872 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_872 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_873 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h369 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_873 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_873 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_874 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_874 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_874 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_875 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_875 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_875 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_876 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_876 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_876 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_877 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_877 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_877 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_878 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_878 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_878 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_879 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h36f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_879 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_879 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_880 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h370 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_880 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_880 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_881 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h371 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_881 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_881 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_882 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h372 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_882 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_882 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_883 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h373 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_883 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_883 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_884 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h374 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_884 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_884 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_885 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h375 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_885 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_885 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_886 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h376 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_886 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_886 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_887 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h377 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_887 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_887 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_888 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h378 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_888 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_888 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_889 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h379 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_889 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_889 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_890 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_890 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_890 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_891 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_891 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_891 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_892 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_892 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_892 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_893 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_893 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_893 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_894 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_894 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_894 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_895 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h37f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_895 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_895 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_896 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h380 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_896 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_896 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_897 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h381 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_897 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_897 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_898 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h382 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_898 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_898 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_899 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h383 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_899 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_899 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_900 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h384 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_900 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_900 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_901 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h385 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_901 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_901 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_902 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h386 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_902 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_902 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_903 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h387 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_903 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_903 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_904 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h388 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_904 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_904 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_905 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h389 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_905 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_905 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_906 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_906 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_906 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_907 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_907 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_907 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_908 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_908 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_908 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_909 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_909 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_909 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_910 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_910 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_910 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_911 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h38f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_911 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_911 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_912 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h390 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_912 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_912 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_913 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h391 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_913 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_913 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_914 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h392 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_914 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_914 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_915 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h393 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_915 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_915 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_916 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h394 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_916 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_916 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_917 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h395 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_917 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_917 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_918 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h396 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_918 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_918 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_919 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h397 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_919 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_919 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_920 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h398 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_920 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_920 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_921 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h399 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_921 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_921 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_922 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_922 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_922 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_923 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_923 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_923 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_924 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_924 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_924 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_925 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_925 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_925 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_926 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_926 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_926 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_927 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h39f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_927 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_927 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_928 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_928 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_928 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_929 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_929 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_929 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_930 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_930 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_930 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_931 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_931 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_931 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_932 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_932 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_932 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_933 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_933 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_933 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_934 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_934 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_934 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_935 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_935 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_935 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_936 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_936 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_936 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_937 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_937 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_937 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_938 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_938 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_938 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_939 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_939 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_939 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_940 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_940 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_940 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_941 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_941 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_941 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_942 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_942 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_942 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_943 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_943 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_943 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_944 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_944 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_944 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_945 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_945 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_945 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_946 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_946 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_946 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_947 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_947 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_947 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_948 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_948 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_948 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_949 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_949 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_949 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_950 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_950 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_950 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_951 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_951 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_951 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_952 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_952 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_952 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_953 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_953 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_953 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_954 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_954 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_954 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_955 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_955 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_955 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_956 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_956 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_956 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_957 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_957 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_957 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_958 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_958 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_958 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_959 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_959 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_959 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_960 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_960 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_960 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_961 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_961 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_961 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_962 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_962 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_962 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_963 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_963 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_963 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_964 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_964 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_964 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_965 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_965 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_965 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_966 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_966 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_966 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_967 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_967 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_967 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_968 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_968 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_968 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_969 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_969 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_969 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_970 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_970 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_970 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_971 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_971 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_971 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_972 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_972 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_972 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_973 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_973 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_973 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_974 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_974 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_974 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_975 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_975 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_975 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_976 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_976 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_976 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_977 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_977 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_977 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_978 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_978 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_978 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_979 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_979 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_979 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_980 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_980 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_980 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_981 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_981 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_981 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_982 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_982 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_982 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_983 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_983 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_983 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_984 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_984 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_984 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_985 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_985 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_985 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_986 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_986 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_986 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_987 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_987 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_987 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_988 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_988 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_988 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_989 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_989 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_989 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_990 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_990 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_990 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_991 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_991 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_991 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_992 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_992 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_992 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_993 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_993 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_993 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_994 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_994 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_994 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_995 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_995 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_995 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_996 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_996 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_996 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_997 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_997 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_997 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_998 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_998 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_998 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_999 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_999 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_999 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1000 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1000 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1000 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1001 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1001 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1001 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1002 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1002 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1002 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1003 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1003 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1003 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1004 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1004 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1004 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1005 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1005 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1005 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1006 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1006 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1006 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1007 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1007 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1007 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1008 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1008 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1008 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1009 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1009 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1009 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1010 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1010 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1010 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1011 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1011 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1011 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1012 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1012 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1012 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1013 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1013 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1013 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1014 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1014 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1014 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1015 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1015 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1015 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1016 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1016 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1016 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1017 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1017 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1017 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1018 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1018 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1018 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1019 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1019 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1019 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1020 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1020 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1020 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1021 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1021 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1021 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1022 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1022 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1022 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1023 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h3ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1023 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1023 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1024 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h400 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1024 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1024 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1025 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h401 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1025 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1025 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1026 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h402 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1026 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1026 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1027 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h403 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1027 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1027 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1028 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h404 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1028 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1028 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1029 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h405 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1029 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1029 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1030 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h406 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1030 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1030 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1031 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h407 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1031 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1031 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1032 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h408 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1032 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1032 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1033 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h409 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1033 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1033 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1034 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1034 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1034 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1035 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1035 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1035 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1036 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1036 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1036 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1037 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1037 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1037 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1038 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1038 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1038 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1039 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h40f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1039 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1039 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1040 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h410 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1040 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1040 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1041 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h411 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1041 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1041 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1042 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h412 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1042 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1042 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1043 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h413 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1043 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1043 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1044 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h414 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1044 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1044 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1045 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h415 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1045 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1045 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1046 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h416 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1046 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1046 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1047 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h417 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1047 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1047 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1048 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h418 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1048 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1048 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1049 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h419 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1049 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1049 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1050 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1050 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1050 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1051 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1051 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1051 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1052 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1052 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1052 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1053 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1053 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1053 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1054 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1054 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1054 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1055 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h41f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1055 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1055 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1056 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h420 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1056 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1056 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1057 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h421 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1057 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1057 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1058 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h422 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1058 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1058 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1059 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h423 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1059 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1059 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1060 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h424 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1060 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1060 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1061 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h425 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1061 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1061 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1062 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h426 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1062 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1062 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1063 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h427 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1063 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1063 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1064 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h428 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1064 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1064 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1065 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h429 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1065 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1065 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1066 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1066 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1066 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1067 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1067 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1067 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1068 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1068 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1068 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1069 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1069 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1069 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1070 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1070 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1070 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1071 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h42f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1071 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1071 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1072 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h430 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1072 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1072 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1073 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h431 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1073 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1073 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1074 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h432 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1074 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1074 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1075 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h433 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1075 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1075 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1076 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h434 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1076 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1076 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1077 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h435 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1077 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1077 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1078 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h436 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1078 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1078 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1079 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h437 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1079 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1079 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1080 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h438 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1080 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1080 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1081 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h439 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1081 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1081 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1082 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1082 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1082 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1083 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1083 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1083 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1084 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1084 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1084 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1085 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1085 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1085 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1086 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1086 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1086 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1087 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h43f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1087 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1087 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1088 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h440 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1088 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1088 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1089 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h441 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1089 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1089 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1090 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h442 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1090 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1090 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1091 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h443 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1091 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1091 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1092 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h444 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1092 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1092 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1093 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h445 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1093 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1093 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1094 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h446 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1094 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1094 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1095 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h447 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1095 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1095 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1096 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h448 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1096 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1096 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1097 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h449 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1097 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1097 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1098 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1098 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1098 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1099 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1099 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1099 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1100 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1100 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1100 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1101 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1101 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1101 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1102 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1102 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1102 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1103 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h44f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1103 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1103 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1104 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h450 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1104 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1104 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1105 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h451 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1105 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1105 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1106 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h452 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1106 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1106 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1107 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h453 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1107 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1107 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1108 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h454 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1108 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1108 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1109 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h455 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1109 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1109 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1110 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h456 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1110 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1110 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1111 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h457 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1111 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1111 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1112 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h458 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1112 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1112 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1113 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h459 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1113 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1113 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1114 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1114 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1114 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1115 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1115 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1115 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1116 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1116 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1116 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1117 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1117 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1117 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1118 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1118 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1118 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1119 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h45f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1119 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1119 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1120 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h460 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1120 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1120 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1121 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h461 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1121 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1121 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1122 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h462 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1122 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1122 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1123 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h463 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1123 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1123 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1124 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h464 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1124 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1124 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1125 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h465 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1125 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1125 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1126 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h466 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1126 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1126 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1127 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h467 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1127 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1127 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1128 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h468 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1128 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1128 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1129 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h469 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1129 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1129 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1130 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1130 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1130 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1131 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1131 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1131 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1132 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1132 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1132 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1133 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1133 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1133 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1134 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1134 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1134 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1135 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h46f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1135 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1135 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1136 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h470 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1136 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1136 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1137 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h471 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1137 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1137 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1138 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h472 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1138 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1138 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1139 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h473 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1139 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1139 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1140 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h474 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1140 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1140 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1141 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h475 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1141 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1141 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1142 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h476 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1142 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1142 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1143 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h477 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1143 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1143 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1144 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h478 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1144 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1144 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1145 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h479 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1145 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1145 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1146 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1146 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1146 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1147 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1147 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1147 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1148 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1148 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1148 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1149 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1149 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1149 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1150 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1150 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1150 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1151 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h47f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1151 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1151 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1152 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h480 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1152 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1152 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1153 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h481 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1153 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1153 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1154 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h482 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1154 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1154 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1155 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h483 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1155 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1155 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1156 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h484 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1156 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1156 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1157 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h485 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1157 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1157 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1158 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h486 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1158 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1158 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1159 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h487 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1159 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1159 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1160 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h488 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1160 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1160 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1161 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h489 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1161 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1161 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1162 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1162 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1162 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1163 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1163 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1163 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1164 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1164 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1164 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1165 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1165 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1165 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1166 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1166 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1166 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1167 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h48f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1167 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1167 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1168 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h490 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1168 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1168 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1169 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h491 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1169 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1169 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1170 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h492 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1170 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1170 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1171 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h493 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1171 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1171 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1172 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h494 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1172 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1172 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1173 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h495 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1173 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1173 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1174 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h496 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1174 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1174 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1175 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h497 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1175 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1175 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1176 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h498 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1176 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1176 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1177 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h499 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1177 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1177 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1178 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1178 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1178 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1179 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1179 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1179 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1180 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1180 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1180 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1181 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1181 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1181 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1182 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1182 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1182 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1183 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h49f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1183 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1183 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1184 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1184 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1184 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1185 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1185 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1185 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1186 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1186 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1186 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1187 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1187 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1187 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1188 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1188 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1188 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1189 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1189 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1189 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1190 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1190 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1190 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1191 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1191 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1191 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1192 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1192 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1192 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1193 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1193 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1193 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1194 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1194 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1194 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1195 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1195 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1195 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1196 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1196 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1196 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1197 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1197 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1197 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1198 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1198 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1198 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1199 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1199 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1199 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1200 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1200 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1200 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1201 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1201 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1201 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1202 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1202 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1202 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1203 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1203 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1203 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1204 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1204 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1204 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1205 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1205 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1205 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1206 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1206 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1206 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1207 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1207 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1207 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1208 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1208 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1208 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1209 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1209 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1209 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1210 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1210 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1210 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1211 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1211 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1211 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1212 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1212 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1212 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1213 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1213 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1213 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1214 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1214 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1214 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1215 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1215 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1215 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1216 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1216 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1216 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1217 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1217 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1217 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1218 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1218 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1218 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1219 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1219 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1219 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1220 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1220 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1220 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1221 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1221 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1221 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1222 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1222 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1222 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1223 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1223 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1223 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1224 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1224 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1224 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1225 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1225 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1225 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1226 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1226 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1226 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1227 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1227 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1227 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1228 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1228 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1228 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1229 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1229 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1229 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1230 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1230 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1230 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1231 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1231 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1231 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1232 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1232 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1232 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1233 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1233 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1233 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1234 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1234 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1234 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1235 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1235 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1235 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1236 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1236 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1236 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1237 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1237 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1237 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1238 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1238 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1238 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1239 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1239 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1239 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1240 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1240 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1240 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1241 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1241 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1241 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1242 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1242 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1242 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1243 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1243 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1243 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1244 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1244 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1244 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1245 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1245 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1245 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1246 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1246 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1246 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1247 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1247 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1247 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1248 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1248 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1248 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1249 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1249 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1249 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1250 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1250 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1250 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1251 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1251 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1251 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1252 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1252 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1252 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1253 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1253 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1253 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1254 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1254 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1254 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1255 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1255 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1255 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1256 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1256 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1256 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1257 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1257 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1257 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1258 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1258 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1258 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1259 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1259 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1259 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1260 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1260 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1260 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1261 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1261 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1261 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1262 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1262 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1262 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1263 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1263 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1263 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1264 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1264 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1264 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1265 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1265 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1265 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1266 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1266 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1266 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1267 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1267 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1267 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1268 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1268 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1268 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1269 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1269 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1269 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1270 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1270 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1270 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1271 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1271 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1271 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1272 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1272 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1272 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1273 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1273 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1273 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1274 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1274 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1274 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1275 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1275 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1275 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1276 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1276 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1276 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1277 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1277 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1277 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1278 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1278 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1278 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1279 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h4ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1279 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1279 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1280 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h500 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1280 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1280 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1281 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h501 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1281 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1281 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1282 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h502 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1282 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1282 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1283 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h503 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1283 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1283 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1284 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h504 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1284 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1284 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1285 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h505 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1285 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1285 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1286 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h506 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1286 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1286 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1287 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h507 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1287 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1287 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1288 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h508 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1288 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1288 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1289 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h509 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1289 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1289 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1290 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1290 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1290 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1291 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1291 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1291 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1292 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1292 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1292 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1293 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1293 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1293 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1294 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1294 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1294 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1295 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h50f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1295 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1295 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1296 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h510 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1296 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1296 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1297 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h511 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1297 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1297 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1298 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h512 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1298 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1298 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1299 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h513 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1299 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1299 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1300 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h514 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1300 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1300 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1301 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h515 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1301 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1301 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1302 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h516 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1302 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1302 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1303 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h517 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1303 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1303 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1304 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h518 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1304 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1304 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1305 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h519 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1305 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1305 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1306 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1306 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1306 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1307 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1307 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1307 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1308 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1308 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1308 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1309 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1309 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1309 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1310 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1310 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1310 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1311 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h51f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1311 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1311 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1312 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h520 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1312 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1312 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1313 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h521 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1313 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1313 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1314 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h522 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1314 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1314 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1315 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h523 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1315 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1315 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1316 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h524 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1316 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1316 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1317 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h525 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1317 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1317 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1318 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h526 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1318 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1318 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1319 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h527 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1319 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1319 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1320 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h528 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1320 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1320 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1321 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h529 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1321 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1321 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1322 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1322 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1322 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1323 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1323 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1323 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1324 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1324 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1324 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1325 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1325 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1325 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1326 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1326 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1326 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1327 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h52f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1327 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1327 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1328 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h530 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1328 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1328 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1329 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h531 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1329 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1329 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1330 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h532 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1330 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1330 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1331 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h533 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1331 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1331 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1332 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h534 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1332 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1332 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1333 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h535 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1333 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1333 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1334 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h536 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1334 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1334 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1335 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h537 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1335 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1335 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1336 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h538 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1336 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1336 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1337 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h539 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1337 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1337 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1338 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1338 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1338 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1339 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1339 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1339 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1340 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1340 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1340 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1341 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1341 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1341 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1342 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1342 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1342 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1343 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h53f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1343 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1343 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1344 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h540 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1344 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1344 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1345 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h541 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1345 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1345 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1346 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h542 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1346 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1346 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1347 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h543 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1347 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1347 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1348 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h544 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1348 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1348 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1349 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h545 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1349 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1349 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1350 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h546 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1350 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1350 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1351 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h547 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1351 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1351 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1352 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h548 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1352 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1352 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1353 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h549 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1353 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1353 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1354 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1354 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1354 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1355 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1355 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1355 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1356 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1356 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1356 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1357 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1357 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1357 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1358 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1358 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1358 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1359 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h54f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1359 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1359 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1360 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h550 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1360 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1360 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1361 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h551 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1361 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1361 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1362 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h552 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1362 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1362 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1363 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h553 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1363 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1363 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1364 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h554 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1364 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1364 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1365 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h555 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1365 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1365 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1366 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h556 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1366 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1366 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1367 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h557 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1367 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1367 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1368 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h558 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1368 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1368 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1369 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h559 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1369 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1369 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1370 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1370 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1370 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1371 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1371 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1371 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1372 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1372 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1372 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1373 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1373 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1373 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1374 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1374 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1374 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1375 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h55f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1375 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1375 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1376 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h560 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1376 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1376 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1377 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h561 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1377 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1377 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1378 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h562 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1378 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1378 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1379 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h563 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1379 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1379 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1380 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h564 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1380 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1380 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1381 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h565 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1381 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1381 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1382 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h566 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1382 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1382 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1383 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h567 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1383 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1383 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1384 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h568 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1384 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1384 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1385 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h569 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1385 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1385 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1386 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1386 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1386 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1387 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1387 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1387 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1388 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1388 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1388 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1389 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1389 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1389 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1390 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1390 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1390 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1391 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h56f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1391 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1391 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1392 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h570 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1392 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1392 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1393 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h571 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1393 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1393 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1394 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h572 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1394 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1394 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1395 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h573 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1395 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1395 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1396 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h574 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1396 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1396 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1397 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h575 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1397 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1397 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1398 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h576 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1398 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1398 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1399 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h577 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1399 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1399 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1400 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h578 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1400 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1400 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1401 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h579 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1401 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1401 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1402 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1402 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1402 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1403 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1403 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1403 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1404 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1404 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1404 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1405 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1405 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1405 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1406 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1406 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1406 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1407 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h57f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1407 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1407 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1408 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h580 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1408 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1408 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1409 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h581 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1409 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1409 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1410 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h582 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1410 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1410 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1411 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h583 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1411 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1411 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1412 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h584 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1412 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1412 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1413 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h585 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1413 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1413 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1414 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h586 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1414 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1414 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1415 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h587 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1415 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1415 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1416 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h588 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1416 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1416 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1417 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h589 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1417 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1417 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1418 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1418 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1418 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1419 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1419 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1419 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1420 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1420 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1420 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1421 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1421 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1421 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1422 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1422 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1422 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1423 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h58f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1423 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1423 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1424 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h590 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1424 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1424 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1425 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h591 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1425 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1425 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1426 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h592 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1426 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1426 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1427 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h593 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1427 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1427 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1428 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h594 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1428 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1428 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1429 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h595 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1429 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1429 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1430 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h596 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1430 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1430 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1431 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h597 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1431 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1431 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1432 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h598 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1432 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1432 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1433 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h599 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1433 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1433 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1434 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1434 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1434 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1435 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1435 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1435 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1436 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1436 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1436 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1437 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1437 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1437 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1438 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1438 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1438 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1439 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h59f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1439 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1439 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1440 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1440 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1440 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1441 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1441 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1441 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1442 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1442 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1442 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1443 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1443 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1443 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1444 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1444 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1444 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1445 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1445 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1445 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1446 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1446 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1446 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1447 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1447 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1447 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1448 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1448 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1448 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1449 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1449 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1449 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1450 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1450 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1450 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1451 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1451 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1451 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1452 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1452 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1452 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1453 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1453 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1453 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1454 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1454 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1454 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1455 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1455 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1455 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1456 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1456 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1456 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1457 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1457 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1457 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1458 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1458 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1458 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1459 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1459 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1459 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1460 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1460 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1460 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1461 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1461 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1461 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1462 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1462 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1462 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1463 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1463 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1463 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1464 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1464 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1464 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1465 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1465 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1465 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1466 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1466 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1466 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1467 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1467 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1467 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1468 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1468 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1468 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1469 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1469 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1469 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1470 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1470 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1470 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1471 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1471 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1471 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1472 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1472 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1472 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1473 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1473 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1473 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1474 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1474 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1474 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1475 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1475 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1475 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1476 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1476 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1476 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1477 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1477 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1477 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1478 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1478 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1478 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1479 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1479 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1479 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1480 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1480 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1480 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1481 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1481 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1481 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1482 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1482 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1482 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1483 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1483 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1483 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1484 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1484 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1484 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1485 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1485 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1485 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1486 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1486 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1486 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1487 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1487 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1487 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1488 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1488 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1488 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1489 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1489 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1489 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1490 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1490 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1490 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1491 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1491 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1491 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1492 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1492 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1492 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1493 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1493 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1493 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1494 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1494 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1494 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1495 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1495 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1495 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1496 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1496 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1496 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1497 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1497 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1497 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1498 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1498 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1498 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1499 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1499 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1499 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1500 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1500 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1500 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1501 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1501 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1501 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1502 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1502 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1502 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1503 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1503 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1503 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1504 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1504 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1504 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1505 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1505 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1505 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1506 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1506 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1506 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1507 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1507 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1507 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1508 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1508 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1508 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1509 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1509 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1509 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1510 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1510 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1510 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1511 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1511 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1511 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1512 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1512 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1512 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1513 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1513 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1513 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1514 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1514 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1514 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1515 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1515 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1515 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1516 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1516 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1516 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1517 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1517 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1517 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1518 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1518 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1518 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1519 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1519 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1519 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1520 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1520 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1520 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1521 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1521 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1521 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1522 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1522 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1522 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1523 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1523 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1523 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1524 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1524 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1524 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1525 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1525 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1525 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1526 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1526 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1526 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1527 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1527 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1527 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1528 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1528 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1528 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1529 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1529 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1529 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1530 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1530 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1530 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1531 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1531 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1531 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1532 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1532 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1532 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1533 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1533 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1533 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1534 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1534 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1534 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1535 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h5ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1535 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1535 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1536 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h600 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1536 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1536 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1537 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h601 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1537 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1537 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1538 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h602 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1538 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1538 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1539 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h603 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1539 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1539 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1540 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h604 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1540 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1540 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1541 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h605 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1541 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1541 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1542 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h606 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1542 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1542 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1543 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h607 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1543 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1543 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1544 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h608 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1544 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1544 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1545 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h609 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1545 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1545 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1546 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1546 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1546 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1547 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1547 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1547 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1548 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1548 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1548 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1549 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1549 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1549 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1550 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1550 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1550 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1551 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h60f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1551 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1551 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1552 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h610 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1552 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1552 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1553 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h611 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1553 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1553 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1554 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h612 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1554 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1554 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1555 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h613 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1555 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1555 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1556 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h614 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1556 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1556 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1557 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h615 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1557 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1557 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1558 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h616 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1558 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1558 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1559 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h617 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1559 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1559 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1560 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h618 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1560 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1560 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1561 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h619 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1561 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1561 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1562 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1562 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1562 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1563 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1563 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1563 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1564 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1564 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1564 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1565 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1565 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1565 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1566 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1566 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1566 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1567 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h61f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1567 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1567 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1568 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h620 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1568 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1568 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1569 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h621 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1569 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1569 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1570 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h622 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1570 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1570 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1571 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h623 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1571 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1571 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1572 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h624 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1572 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1572 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1573 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h625 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1573 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1573 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1574 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h626 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1574 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1574 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1575 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h627 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1575 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1575 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1576 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h628 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1576 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1576 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1577 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h629 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1577 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1577 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1578 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1578 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1578 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1579 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1579 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1579 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1580 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1580 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1580 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1581 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1581 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1581 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1582 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1582 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1582 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1583 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h62f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1583 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1583 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1584 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h630 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1584 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1584 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1585 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h631 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1585 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1585 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1586 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h632 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1586 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1586 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1587 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h633 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1587 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1587 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1588 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h634 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1588 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1588 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1589 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h635 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1589 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1589 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1590 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h636 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1590 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1590 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1591 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h637 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1591 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1591 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1592 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h638 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1592 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1592 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1593 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h639 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1593 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1593 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1594 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1594 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1594 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1595 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1595 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1595 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1596 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1596 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1596 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1597 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1597 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1597 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1598 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1598 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1598 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1599 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h63f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1599 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1599 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1600 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h640 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1600 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1600 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1601 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h641 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1601 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1601 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1602 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h642 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1602 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1602 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1603 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h643 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1603 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1603 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1604 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h644 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1604 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1604 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1605 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h645 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1605 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1605 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1606 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h646 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1606 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1606 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1607 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h647 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1607 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1607 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1608 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h648 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1608 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1608 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1609 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h649 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1609 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1609 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1610 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1610 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1610 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1611 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1611 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1611 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1612 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1612 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1612 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1613 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1613 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1613 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1614 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1614 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1614 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1615 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h64f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1615 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1615 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1616 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h650 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1616 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1616 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1617 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h651 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1617 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1617 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1618 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h652 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1618 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1618 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1619 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h653 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1619 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1619 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1620 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h654 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1620 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1620 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1621 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h655 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1621 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1621 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1622 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h656 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1622 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1622 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1623 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h657 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1623 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1623 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1624 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h658 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1624 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1624 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1625 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h659 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1625 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1625 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1626 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1626 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1626 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1627 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1627 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1627 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1628 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1628 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1628 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1629 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1629 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1629 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1630 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1630 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1630 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1631 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h65f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1631 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1631 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1632 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h660 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1632 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1632 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1633 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h661 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1633 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1633 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1634 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h662 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1634 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1634 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1635 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h663 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1635 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1635 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1636 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h664 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1636 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1636 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1637 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h665 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1637 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1637 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1638 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h666 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1638 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1638 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1639 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h667 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1639 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1639 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1640 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h668 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1640 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1640 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1641 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h669 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1641 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1641 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1642 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1642 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1642 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1643 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1643 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1643 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1644 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1644 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1644 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1645 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1645 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1645 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1646 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1646 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1646 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1647 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h66f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1647 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1647 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1648 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h670 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1648 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1648 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1649 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h671 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1649 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1649 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1650 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h672 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1650 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1650 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1651 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h673 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1651 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1651 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1652 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h674 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1652 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1652 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1653 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h675 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1653 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1653 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1654 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h676 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1654 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1654 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1655 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h677 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1655 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1655 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1656 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h678 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1656 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1656 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1657 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h679 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1657 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1657 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1658 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1658 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1658 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1659 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1659 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1659 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1660 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1660 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1660 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1661 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1661 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1661 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1662 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1662 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1662 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1663 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h67f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1663 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1663 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1664 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h680 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1664 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1664 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1665 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h681 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1665 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1665 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1666 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h682 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1666 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1666 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1667 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h683 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1667 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1667 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1668 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h684 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1668 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1668 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1669 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h685 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1669 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1669 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1670 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h686 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1670 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1670 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1671 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h687 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1671 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1671 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1672 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h688 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1672 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1672 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1673 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h689 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1673 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1673 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1674 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1674 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1674 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1675 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1675 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1675 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1676 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1676 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1676 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1677 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1677 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1677 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1678 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1678 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1678 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1679 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h68f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1679 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1679 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1680 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h690 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1680 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1680 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1681 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h691 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1681 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1681 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1682 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h692 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1682 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1682 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1683 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h693 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1683 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1683 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1684 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h694 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1684 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1684 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1685 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h695 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1685 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1685 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1686 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h696 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1686 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1686 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1687 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h697 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1687 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1687 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1688 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h698 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1688 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1688 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1689 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h699 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1689 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1689 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1690 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1690 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1690 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1691 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1691 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1691 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1692 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1692 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1692 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1693 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1693 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1693 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1694 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1694 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1694 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1695 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h69f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1695 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1695 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1696 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1696 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1696 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1697 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1697 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1697 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1698 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1698 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1698 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1699 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1699 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1699 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1700 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1700 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1700 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1701 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1701 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1701 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1702 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1702 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1702 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1703 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1703 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1703 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1704 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1704 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1704 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1705 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1705 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1705 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1706 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1706 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1706 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1707 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1707 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1707 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1708 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1708 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1708 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1709 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1709 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1709 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1710 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1710 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1710 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1711 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1711 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1711 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1712 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1712 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1712 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1713 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1713 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1713 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1714 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1714 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1714 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1715 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1715 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1715 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1716 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1716 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1716 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1717 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1717 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1717 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1718 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1718 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1718 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1719 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1719 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1719 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1720 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1720 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1720 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1721 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1721 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1721 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1722 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1722 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1722 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1723 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1723 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1723 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1724 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1724 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1724 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1725 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1725 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1725 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1726 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1726 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1726 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1727 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1727 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1727 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1728 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1728 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1728 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1729 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1729 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1729 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1730 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1730 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1730 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1731 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1731 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1731 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1732 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1732 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1732 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1733 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1733 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1733 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1734 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1734 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1734 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1735 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1735 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1735 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1736 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1736 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1736 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1737 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1737 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1737 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1738 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1738 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1738 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1739 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1739 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1739 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1740 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1740 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1740 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1741 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1741 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1741 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1742 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1742 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1742 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1743 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1743 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1743 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1744 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1744 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1744 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1745 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1745 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1745 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1746 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1746 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1746 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1747 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1747 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1747 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1748 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1748 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1748 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1749 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1749 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1749 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1750 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1750 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1750 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1751 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1751 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1751 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1752 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1752 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1752 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1753 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1753 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1753 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1754 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1754 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1754 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1755 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1755 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1755 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1756 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1756 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1756 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1757 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1757 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1757 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1758 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1758 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1758 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1759 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1759 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1759 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1760 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1760 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1760 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1761 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1761 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1761 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1762 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1762 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1762 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1763 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1763 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1763 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1764 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1764 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1764 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1765 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1765 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1765 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1766 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1766 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1766 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1767 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1767 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1767 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1768 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1768 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1768 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1769 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1769 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1769 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1770 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1770 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1770 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1771 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1771 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1771 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1772 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1772 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1772 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1773 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1773 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1773 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1774 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1774 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1774 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1775 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1775 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1775 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1776 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1776 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1776 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1777 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1777 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1777 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1778 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1778 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1778 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1779 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1779 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1779 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1780 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1780 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1780 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1781 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1781 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1781 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1782 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1782 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1782 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1783 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1783 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1783 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1784 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1784 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1784 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1785 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1785 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1785 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1786 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1786 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1786 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1787 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1787 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1787 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1788 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1788 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1788 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1789 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1789 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1789 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1790 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1790 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1790 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1791 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h6ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1791 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1791 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1792 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h700 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1792 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1792 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1793 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h701 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1793 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1793 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1794 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h702 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1794 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1794 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1795 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h703 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1795 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1795 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1796 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h704 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1796 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1796 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1797 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h705 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1797 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1797 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1798 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h706 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1798 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1798 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1799 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h707 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1799 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1799 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1800 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h708 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1800 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1800 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1801 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h709 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1801 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1801 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1802 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1802 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1802 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1803 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1803 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1803 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1804 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1804 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1804 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1805 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1805 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1805 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1806 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1806 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1806 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1807 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h70f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1807 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1807 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1808 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h710 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1808 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1808 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1809 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h711 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1809 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1809 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1810 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h712 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1810 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1810 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1811 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h713 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1811 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1811 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1812 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h714 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1812 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1812 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1813 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h715 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1813 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1813 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1814 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h716 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1814 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1814 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1815 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h717 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1815 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1815 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1816 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h718 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1816 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1816 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1817 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h719 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1817 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1817 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1818 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1818 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1818 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1819 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1819 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1819 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1820 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1820 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1820 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1821 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1821 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1821 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1822 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1822 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1822 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1823 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h71f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1823 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1823 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1824 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h720 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1824 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1824 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1825 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h721 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1825 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1825 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1826 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h722 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1826 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1826 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1827 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h723 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1827 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1827 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1828 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h724 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1828 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1828 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1829 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h725 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1829 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1829 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1830 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h726 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1830 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1830 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1831 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h727 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1831 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1831 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1832 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h728 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1832 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1832 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1833 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h729 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1833 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1833 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1834 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1834 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1834 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1835 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1835 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1835 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1836 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1836 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1836 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1837 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1837 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1837 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1838 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1838 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1838 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1839 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h72f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1839 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1839 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1840 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h730 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1840 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1840 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1841 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h731 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1841 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1841 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1842 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h732 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1842 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1842 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1843 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h733 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1843 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1843 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1844 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h734 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1844 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1844 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1845 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h735 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1845 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1845 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1846 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h736 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1846 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1846 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1847 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h737 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1847 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1847 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1848 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h738 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1848 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1848 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1849 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h739 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1849 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1849 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1850 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1850 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1850 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1851 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1851 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1851 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1852 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1852 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1852 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1853 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1853 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1853 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1854 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1854 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1854 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1855 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h73f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1855 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1855 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1856 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h740 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1856 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1856 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1857 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h741 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1857 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1857 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1858 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h742 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1858 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1858 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1859 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h743 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1859 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1859 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1860 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h744 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1860 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1860 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1861 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h745 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1861 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1861 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1862 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h746 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1862 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1862 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1863 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h747 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1863 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1863 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1864 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h748 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1864 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1864 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1865 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h749 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1865 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1865 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1866 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1866 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1866 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1867 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1867 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1867 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1868 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1868 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1868 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1869 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1869 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1869 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1870 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1870 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1870 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1871 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h74f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1871 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1871 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1872 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h750 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1872 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1872 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1873 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h751 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1873 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1873 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1874 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h752 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1874 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1874 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1875 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h753 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1875 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1875 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1876 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h754 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1876 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1876 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1877 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h755 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1877 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1877 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1878 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h756 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1878 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1878 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1879 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h757 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1879 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1879 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1880 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h758 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1880 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1880 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1881 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h759 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1881 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1881 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1882 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1882 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1882 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1883 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1883 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1883 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1884 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1884 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1884 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1885 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1885 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1885 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1886 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1886 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1886 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1887 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h75f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1887 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1887 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1888 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h760 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1888 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1888 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1889 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h761 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1889 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1889 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1890 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h762 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1890 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1890 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1891 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h763 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1891 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1891 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1892 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h764 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1892 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1892 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1893 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h765 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1893 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1893 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1894 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h766 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1894 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1894 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1895 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h767 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1895 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1895 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1896 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h768 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1896 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1896 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1897 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h769 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1897 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1897 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1898 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1898 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1898 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1899 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1899 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1899 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1900 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1900 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1900 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1901 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1901 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1901 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1902 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1902 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1902 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1903 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h76f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1903 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1903 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1904 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h770 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1904 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1904 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1905 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h771 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1905 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1905 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1906 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h772 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1906 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1906 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1907 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h773 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1907 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1907 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1908 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h774 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1908 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1908 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1909 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h775 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1909 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1909 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1910 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h776 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1910 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1910 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1911 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h777 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1911 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1911 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1912 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h778 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1912 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1912 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1913 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h779 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1913 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1913 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1914 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1914 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1914 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1915 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1915 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1915 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1916 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1916 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1916 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1917 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1917 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1917 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1918 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1918 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1918 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1919 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h77f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1919 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1919 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1920 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h780 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1920 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1920 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1921 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h781 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1921 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1921 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1922 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h782 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1922 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1922 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1923 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h783 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1923 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1923 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1924 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h784 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1924 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1924 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1925 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h785 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1925 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1925 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1926 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h786 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1926 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1926 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1927 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h787 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1927 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1927 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1928 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h788 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1928 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1928 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1929 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h789 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1929 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1929 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1930 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1930 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1930 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1931 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1931 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1931 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1932 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1932 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1932 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1933 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1933 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1933 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1934 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1934 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1934 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1935 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h78f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1935 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1935 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1936 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h790 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1936 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1936 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1937 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h791 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1937 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1937 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1938 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h792 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1938 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1938 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1939 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h793 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1939 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1939 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1940 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h794 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1940 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1940 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1941 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h795 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1941 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1941 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1942 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h796 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1942 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1942 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1943 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h797 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1943 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1943 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1944 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h798 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1944 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1944 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1945 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h799 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1945 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1945 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1946 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1946 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1946 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1947 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1947 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1947 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1948 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1948 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1948 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1949 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1949 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1949 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1950 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1950 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1950 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1951 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h79f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1951 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1951 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1952 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1952 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1952 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1953 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1953 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1953 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1954 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1954 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1954 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1955 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1955 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1955 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1956 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1956 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1956 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1957 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1957 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1957 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1958 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1958 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1958 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1959 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1959 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1959 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1960 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1960 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1960 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1961 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1961 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1961 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1962 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1962 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1962 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1963 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1963 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1963 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1964 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1964 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1964 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1965 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1965 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1965 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1966 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1966 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1966 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1967 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1967 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1967 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1968 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1968 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1968 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1969 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1969 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1969 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1970 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1970 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1970 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1971 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1971 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1971 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1972 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1972 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1972 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1973 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1973 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1973 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1974 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1974 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1974 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1975 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1975 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1975 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1976 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1976 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1976 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1977 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1977 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1977 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1978 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1978 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1978 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1979 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1979 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1979 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1980 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1980 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1980 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1981 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1981 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1981 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1982 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1982 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1982 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1983 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1983 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1983 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1984 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1984 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1984 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1985 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1985 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1985 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1986 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1986 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1986 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1987 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1987 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1987 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1988 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1988 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1988 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1989 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1989 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1989 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1990 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1990 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1990 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1991 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1991 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1991 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1992 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1992 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1992 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1993 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1993 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1993 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1994 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1994 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1994 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1995 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1995 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1995 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1996 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1996 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1996 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1997 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1997 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1997 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1998 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1998 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1998 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_1999 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_1999 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_1999 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2000 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2000 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2000 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2001 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2001 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2001 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2002 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2002 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2002 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2003 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2003 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2003 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2004 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2004 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2004 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2005 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2005 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2005 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2006 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2006 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2006 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2007 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2007 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2007 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2008 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2008 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2008 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2009 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2009 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2009 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2010 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2010 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2010 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2011 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2011 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2011 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2012 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2012 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2012 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2013 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2013 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2013 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2014 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2014 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2014 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2015 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2015 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2015 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2016 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2016 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2016 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2017 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2017 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2017 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2018 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2018 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2018 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2019 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2019 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2019 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2020 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2020 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2020 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2021 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2021 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2021 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2022 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2022 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2022 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2023 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2023 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2023 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2024 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2024 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2024 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2025 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2025 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2025 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2026 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2026 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2026 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2027 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2027 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2027 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2028 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2028 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2028 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2029 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2029 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2029 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2030 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2030 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2030 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2031 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2031 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2031 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2032 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2032 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2032 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2033 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2033 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2033 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2034 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2034 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2034 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2035 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2035 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2035 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2036 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2036 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2036 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2037 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2037 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2037 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2038 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2038 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2038 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2039 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2039 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2039 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2040 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2040 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2040 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2041 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2041 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2041 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2042 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2042 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2042 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2043 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2043 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2043 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2044 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2044 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2044 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2045 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2045 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2045 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2046 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2046 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2046 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2047 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h7ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2047 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2047 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2048 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h800 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2048 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2048 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2049 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h801 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2049 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2049 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2050 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h802 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2050 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2050 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2051 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h803 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2051 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2051 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2052 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h804 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2052 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2052 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2053 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h805 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2053 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2053 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2054 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h806 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2054 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2054 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2055 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h807 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2055 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2055 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2056 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h808 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2056 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2056 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2057 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h809 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2057 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2057 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2058 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2058 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2058 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2059 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2059 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2059 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2060 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2060 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2060 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2061 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2061 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2061 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2062 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2062 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2062 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2063 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h80f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2063 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2063 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2064 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h810 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2064 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2064 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2065 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h811 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2065 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2065 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2066 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h812 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2066 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2066 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2067 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h813 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2067 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2067 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2068 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h814 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2068 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2068 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2069 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h815 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2069 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2069 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2070 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h816 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2070 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2070 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2071 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h817 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2071 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2071 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2072 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h818 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2072 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2072 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2073 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h819 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2073 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2073 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2074 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2074 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2074 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2075 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2075 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2075 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2076 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2076 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2076 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2077 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2077 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2077 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2078 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2078 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2078 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2079 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h81f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2079 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2079 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2080 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h820 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2080 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2080 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2081 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h821 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2081 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2081 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2082 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h822 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2082 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2082 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2083 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h823 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2083 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2083 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2084 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h824 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2084 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2084 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2085 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h825 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2085 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2085 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2086 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h826 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2086 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2086 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2087 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h827 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2087 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2087 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2088 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h828 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2088 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2088 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2089 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h829 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2089 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2089 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2090 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2090 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2090 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2091 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2091 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2091 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2092 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2092 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2092 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2093 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2093 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2093 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2094 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2094 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2094 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2095 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h82f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2095 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2095 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2096 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h830 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2096 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2096 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2097 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h831 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2097 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2097 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2098 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h832 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2098 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2098 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2099 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h833 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2099 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2099 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2100 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h834 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2100 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2100 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2101 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h835 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2101 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2101 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2102 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h836 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2102 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2102 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2103 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h837 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2103 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2103 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2104 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h838 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2104 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2104 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2105 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h839 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2105 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2105 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2106 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2106 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2106 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2107 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2107 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2107 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2108 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2108 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2108 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2109 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2109 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2109 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2110 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2110 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2110 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2111 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h83f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2111 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2111 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2112 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h840 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2112 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2112 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2113 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h841 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2113 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2113 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2114 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h842 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2114 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2114 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2115 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h843 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2115 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2115 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2116 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h844 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2116 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2116 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2117 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h845 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2117 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2117 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2118 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h846 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2118 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2118 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2119 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h847 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2119 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2119 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2120 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h848 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2120 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2120 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2121 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h849 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2121 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2121 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2122 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2122 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2122 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2123 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2123 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2123 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2124 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2124 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2124 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2125 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2125 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2125 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2126 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2126 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2126 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2127 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h84f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2127 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2127 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2128 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h850 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2128 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2128 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2129 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h851 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2129 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2129 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2130 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h852 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2130 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2130 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2131 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h853 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2131 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2131 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2132 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h854 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2132 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2132 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2133 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h855 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2133 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2133 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2134 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h856 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2134 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2134 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2135 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h857 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2135 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2135 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2136 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h858 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2136 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2136 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2137 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h859 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2137 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2137 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2138 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2138 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2138 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2139 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2139 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2139 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2140 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2140 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2140 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2141 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2141 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2141 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2142 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2142 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2142 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2143 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h85f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2143 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2143 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2144 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h860 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2144 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2144 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2145 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h861 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2145 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2145 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2146 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h862 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2146 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2146 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2147 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h863 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2147 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2147 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2148 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h864 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2148 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2148 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2149 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h865 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2149 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2149 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2150 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h866 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2150 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2150 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2151 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h867 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2151 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2151 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2152 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h868 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2152 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2152 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2153 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h869 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2153 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2153 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2154 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2154 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2154 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2155 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2155 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2155 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2156 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2156 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2156 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2157 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2157 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2157 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2158 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2158 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2158 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2159 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h86f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2159 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2159 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2160 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h870 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2160 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2160 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2161 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h871 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2161 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2161 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2162 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h872 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2162 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2162 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2163 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h873 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2163 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2163 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2164 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h874 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2164 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2164 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2165 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h875 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2165 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2165 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2166 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h876 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2166 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2166 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2167 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h877 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2167 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2167 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2168 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h878 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2168 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2168 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2169 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h879 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2169 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2169 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2170 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2170 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2170 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2171 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2171 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2171 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2172 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2172 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2172 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2173 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2173 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2173 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2174 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2174 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2174 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2175 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h87f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2175 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2175 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2176 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h880 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2176 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2176 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2177 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h881 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2177 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2177 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2178 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h882 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2178 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2178 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2179 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h883 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2179 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2179 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2180 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h884 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2180 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2180 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2181 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h885 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2181 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2181 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2182 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h886 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2182 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2182 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2183 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h887 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2183 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2183 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2184 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h888 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2184 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2184 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2185 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h889 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2185 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2185 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2186 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2186 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2186 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2187 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2187 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2187 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2188 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2188 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2188 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2189 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2189 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2189 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2190 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2190 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2190 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2191 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h88f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2191 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2191 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2192 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h890 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2192 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2192 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2193 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h891 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2193 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2193 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2194 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h892 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2194 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2194 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2195 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h893 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2195 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2195 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2196 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h894 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2196 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2196 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2197 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h895 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2197 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2197 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2198 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h896 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2198 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2198 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2199 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h897 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2199 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2199 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2200 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h898 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2200 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2200 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2201 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h899 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2201 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2201 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2202 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2202 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2202 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2203 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2203 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2203 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2204 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2204 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2204 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2205 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2205 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2205 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2206 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2206 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2206 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2207 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h89f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2207 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2207 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2208 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2208 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2208 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2209 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2209 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2209 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2210 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2210 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2210 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2211 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2211 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2211 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2212 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2212 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2212 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2213 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2213 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2213 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2214 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2214 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2214 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2215 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2215 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2215 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2216 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2216 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2216 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2217 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2217 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2217 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2218 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2218 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2218 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2219 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2219 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2219 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2220 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2220 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2220 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2221 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2221 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2221 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2222 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2222 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2222 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2223 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2223 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2223 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2224 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2224 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2224 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2225 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2225 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2225 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2226 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2226 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2226 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2227 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2227 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2227 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2228 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2228 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2228 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2229 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2229 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2229 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2230 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2230 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2230 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2231 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2231 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2231 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2232 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2232 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2232 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2233 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2233 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2233 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2234 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2234 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2234 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2235 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2235 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2235 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2236 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2236 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2236 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2237 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2237 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2237 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2238 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2238 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2238 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2239 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2239 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2239 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2240 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2240 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2240 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2241 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2241 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2241 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2242 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2242 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2242 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2243 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2243 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2243 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2244 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2244 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2244 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2245 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2245 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2245 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2246 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2246 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2246 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2247 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2247 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2247 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2248 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2248 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2248 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2249 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2249 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2249 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2250 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2250 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2250 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2251 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2251 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2251 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2252 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2252 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2252 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2253 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2253 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2253 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2254 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2254 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2254 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2255 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2255 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2255 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2256 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2256 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2256 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2257 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2257 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2257 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2258 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2258 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2258 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2259 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2259 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2259 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2260 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2260 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2260 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2261 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2261 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2261 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2262 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2262 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2262 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2263 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2263 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2263 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2264 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2264 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2264 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2265 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2265 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2265 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2266 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2266 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2266 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2267 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2267 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2267 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2268 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2268 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2268 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2269 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2269 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2269 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2270 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2270 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2270 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2271 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2271 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2271 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2272 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2272 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2272 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2273 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2273 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2273 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2274 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2274 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2274 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2275 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2275 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2275 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2276 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2276 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2276 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2277 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2277 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2277 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2278 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2278 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2278 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2279 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2279 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2279 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2280 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2280 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2280 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2281 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2281 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2281 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2282 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2282 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2282 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2283 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2283 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2283 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2284 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2284 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2284 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2285 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2285 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2285 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2286 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2286 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2286 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2287 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2287 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2287 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2288 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2288 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2288 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2289 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2289 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2289 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2290 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2290 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2290 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2291 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2291 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2291 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2292 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2292 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2292 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2293 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2293 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2293 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2294 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2294 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2294 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2295 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2295 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2295 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2296 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2296 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2296 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2297 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2297 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2297 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2298 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2298 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2298 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2299 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2299 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2299 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2300 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2300 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2300 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2301 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2301 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2301 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2302 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2302 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2302 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2303 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h8ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2303 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2303 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2304 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h900 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2304 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2304 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2305 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h901 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2305 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2305 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2306 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h902 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2306 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2306 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2307 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h903 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2307 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2307 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2308 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h904 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2308 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2308 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2309 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h905 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2309 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2309 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2310 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h906 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2310 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2310 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2311 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h907 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2311 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2311 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2312 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h908 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2312 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2312 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2313 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h909 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2313 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2313 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2314 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2314 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2314 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2315 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2315 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2315 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2316 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2316 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2316 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2317 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2317 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2317 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2318 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2318 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2318 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2319 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h90f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2319 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2319 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2320 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h910 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2320 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2320 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2321 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h911 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2321 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2321 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2322 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h912 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2322 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2322 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2323 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h913 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2323 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2323 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2324 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h914 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2324 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2324 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2325 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h915 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2325 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2325 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2326 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h916 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2326 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2326 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2327 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h917 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2327 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2327 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2328 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h918 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2328 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2328 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2329 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h919 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2329 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2329 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2330 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2330 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2330 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2331 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2331 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2331 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2332 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2332 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2332 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2333 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2333 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2333 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2334 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2334 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2334 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2335 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h91f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2335 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2335 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2336 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h920 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2336 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2336 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2337 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h921 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2337 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2337 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2338 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h922 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2338 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2338 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2339 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h923 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2339 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2339 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2340 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h924 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2340 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2340 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2341 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h925 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2341 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2341 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2342 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h926 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2342 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2342 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2343 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h927 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2343 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2343 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2344 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h928 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2344 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2344 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2345 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h929 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2345 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2345 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2346 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2346 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2346 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2347 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2347 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2347 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2348 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2348 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2348 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2349 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2349 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2349 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2350 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2350 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2350 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2351 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h92f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2351 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2351 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2352 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h930 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2352 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2352 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2353 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h931 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2353 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2353 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2354 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h932 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2354 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2354 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2355 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h933 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2355 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2355 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2356 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h934 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2356 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2356 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2357 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h935 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2357 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2357 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2358 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h936 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2358 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2358 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2359 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h937 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2359 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2359 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2360 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h938 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2360 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2360 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2361 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h939 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2361 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2361 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2362 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2362 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2362 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2363 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2363 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2363 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2364 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2364 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2364 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2365 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2365 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2365 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2366 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2366 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2366 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2367 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h93f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2367 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2367 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2368 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h940 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2368 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2368 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2369 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h941 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2369 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2369 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2370 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h942 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2370 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2370 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2371 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h943 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2371 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2371 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2372 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h944 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2372 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2372 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2373 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h945 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2373 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2373 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2374 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h946 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2374 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2374 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2375 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h947 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2375 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2375 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2376 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h948 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2376 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2376 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2377 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h949 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2377 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2377 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2378 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2378 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2378 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2379 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2379 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2379 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2380 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2380 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2380 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2381 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2381 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2381 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2382 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2382 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2382 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2383 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h94f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2383 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2383 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2384 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h950 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2384 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2384 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2385 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h951 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2385 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2385 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2386 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h952 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2386 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2386 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2387 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h953 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2387 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2387 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2388 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h954 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2388 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2388 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2389 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h955 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2389 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2389 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2390 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h956 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2390 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2390 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2391 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h957 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2391 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2391 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2392 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h958 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2392 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2392 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2393 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h959 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2393 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2393 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2394 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2394 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2394 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2395 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2395 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2395 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2396 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2396 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2396 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2397 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2397 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2397 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2398 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2398 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2398 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2399 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h95f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2399 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2399 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2400 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h960 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2400 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2400 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2401 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h961 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2401 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2401 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2402 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h962 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2402 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2402 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2403 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h963 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2403 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2403 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2404 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h964 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2404 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2404 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2405 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h965 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2405 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2405 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2406 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h966 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2406 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2406 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2407 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h967 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2407 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2407 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2408 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h968 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2408 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2408 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2409 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h969 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2409 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2409 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2410 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2410 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2410 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2411 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2411 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2411 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2412 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2412 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2412 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2413 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2413 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2413 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2414 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2414 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2414 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2415 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h96f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2415 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2415 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2416 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h970 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2416 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2416 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2417 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h971 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2417 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2417 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2418 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h972 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2418 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2418 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2419 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h973 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2419 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2419 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2420 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h974 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2420 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2420 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2421 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h975 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2421 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2421 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2422 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h976 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2422 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2422 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2423 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h977 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2423 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2423 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2424 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h978 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2424 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2424 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2425 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h979 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2425 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2425 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2426 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2426 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2426 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2427 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2427 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2427 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2428 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2428 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2428 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2429 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2429 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2429 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2430 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2430 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2430 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2431 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h97f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2431 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2431 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2432 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h980 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2432 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2432 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2433 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h981 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2433 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2433 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2434 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h982 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2434 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2434 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2435 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h983 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2435 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2435 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2436 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h984 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2436 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2436 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2437 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h985 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2437 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2437 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2438 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h986 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2438 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2438 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2439 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h987 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2439 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2439 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2440 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h988 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2440 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2440 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2441 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h989 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2441 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2441 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2442 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2442 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2442 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2443 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2443 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2443 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2444 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2444 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2444 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2445 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2445 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2445 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2446 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2446 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2446 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2447 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h98f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2447 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2447 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2448 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h990 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2448 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2448 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2449 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h991 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2449 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2449 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2450 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h992 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2450 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2450 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2451 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h993 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2451 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2451 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2452 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h994 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2452 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2452 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2453 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h995 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2453 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2453 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2454 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h996 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2454 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2454 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2455 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h997 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2455 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2455 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2456 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h998 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2456 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2456 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2457 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h999 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2457 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2457 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2458 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2458 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2458 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2459 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2459 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2459 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2460 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2460 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2460 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2461 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2461 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2461 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2462 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2462 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2462 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2463 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h99f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2463 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2463 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2464 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2464 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2464 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2465 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2465 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2465 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2466 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2466 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2466 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2467 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2467 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2467 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2468 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2468 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2468 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2469 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2469 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2469 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2470 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2470 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2470 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2471 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2471 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2471 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2472 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2472 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2472 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2473 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9a9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2473 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2473 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2474 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9aa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2474 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2474 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2475 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2475 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2475 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2476 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2476 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2476 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2477 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2477 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2477 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2478 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2478 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2478 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2479 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9af == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2479 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2479 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2480 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2480 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2480 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2481 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2481 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2481 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2482 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2482 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2482 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2483 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2483 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2483 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2484 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2484 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2484 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2485 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2485 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2485 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2486 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2486 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2486 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2487 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2487 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2487 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2488 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2488 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2488 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2489 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9b9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2489 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2489 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2490 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2490 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2490 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2491 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9bb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2491 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2491 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2492 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9bc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2492 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2492 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2493 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9bd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2493 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2493 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2494 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9be == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2494 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2494 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2495 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9bf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2495 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2495 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2496 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2496 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2496 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2497 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2497 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2497 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2498 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2498 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2498 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2499 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2499 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2499 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2500 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2500 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2500 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2501 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2501 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2501 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2502 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2502 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2502 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2503 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2503 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2503 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2504 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2504 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2504 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2505 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9c9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2505 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2505 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2506 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2506 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2506 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2507 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9cb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2507 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2507 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2508 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9cc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2508 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2508 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2509 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9cd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2509 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2509 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2510 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2510 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2510 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2511 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9cf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2511 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2511 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2512 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2512 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2512 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2513 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2513 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2513 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2514 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2514 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2514 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2515 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2515 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2515 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2516 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2516 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2516 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2517 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2517 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2517 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2518 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2518 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2518 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2519 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2519 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2519 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2520 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2520 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2520 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2521 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9d9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2521 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2521 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2522 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9da == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2522 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2522 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2523 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9db == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2523 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2523 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2524 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9dc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2524 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2524 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2525 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9dd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2525 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2525 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2526 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9de == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2526 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2526 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2527 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9df == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2527 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2527 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2528 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2528 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2528 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2529 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2529 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2529 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2530 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2530 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2530 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2531 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2531 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2531 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2532 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2532 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2532 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2533 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2533 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2533 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2534 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2534 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2534 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2535 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2535 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2535 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2536 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2536 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2536 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2537 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9e9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2537 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2537 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2538 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2538 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2538 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2539 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9eb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2539 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2539 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2540 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2540 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2540 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2541 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2541 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2541 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2542 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2542 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2542 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2543 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2543 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2543 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2544 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2544 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2544 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2545 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2545 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2545 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2546 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2546 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2546 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2547 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2547 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2547 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2548 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2548 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2548 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2549 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2549 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2549 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2550 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2550 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2550 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2551 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2551 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2551 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2552 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2552 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2552 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2553 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9f9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2553 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2553 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2554 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9fa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2554 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2554 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2555 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9fb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2555 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2555 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2556 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9fc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2556 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2556 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2557 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9fd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2557 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2557 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2558 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9fe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2558 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2558 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2559 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'h9ff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2559 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2559 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2560 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2560 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2560 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2561 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2561 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2561 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2562 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2562 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2562 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2563 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2563 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2563 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2564 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2564 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2564 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2565 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2565 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2565 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2566 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2566 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2566 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2567 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2567 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2567 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2568 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2568 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2568 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2569 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2569 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2569 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2570 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2570 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2570 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2571 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2571 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2571 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2572 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2572 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2572 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2573 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2573 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2573 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2574 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2574 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2574 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2575 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2575 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2575 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2576 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2576 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2576 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2577 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2577 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2577 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2578 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2578 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2578 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2579 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2579 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2579 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2580 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2580 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2580 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2581 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2581 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2581 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2582 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2582 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2582 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2583 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2583 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2583 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2584 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2584 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2584 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2585 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2585 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2585 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2586 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2586 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2586 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2587 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2587 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2587 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2588 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2588 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2588 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2589 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2589 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2589 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2590 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2590 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2590 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2591 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2591 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2591 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2592 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2592 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2592 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2593 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2593 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2593 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2594 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2594 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2594 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2595 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2595 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2595 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2596 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2596 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2596 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2597 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2597 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2597 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2598 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2598 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2598 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2599 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2599 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2599 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2600 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2600 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2600 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2601 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2601 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2601 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2602 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2602 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2602 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2603 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2603 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2603 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2604 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2604 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2604 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2605 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2605 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2605 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2606 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2606 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2606 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2607 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2607 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2607 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2608 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2608 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2608 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2609 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2609 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2609 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2610 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2610 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2610 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2611 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2611 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2611 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2612 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2612 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2612 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2613 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2613 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2613 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2614 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2614 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2614 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2615 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2615 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2615 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2616 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2616 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2616 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2617 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2617 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2617 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2618 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2618 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2618 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2619 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2619 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2619 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2620 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2620 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2620 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2621 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2621 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2621 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2622 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2622 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2622 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2623 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2623 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2623 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2624 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2624 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2624 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2625 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2625 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2625 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2626 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2626 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2626 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2627 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2627 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2627 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2628 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2628 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2628 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2629 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2629 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2629 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2630 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2630 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2630 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2631 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2631 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2631 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2632 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2632 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2632 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2633 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2633 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2633 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2634 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2634 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2634 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2635 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2635 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2635 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2636 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2636 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2636 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2637 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2637 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2637 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2638 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2638 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2638 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2639 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2639 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2639 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2640 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2640 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2640 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2641 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2641 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2641 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2642 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2642 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2642 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2643 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2643 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2643 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2644 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2644 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2644 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2645 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2645 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2645 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2646 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2646 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2646 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2647 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2647 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2647 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2648 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2648 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2648 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2649 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2649 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2649 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2650 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2650 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2650 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2651 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2651 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2651 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2652 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2652 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2652 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2653 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2653 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2653 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2654 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2654 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2654 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2655 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2655 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2655 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2656 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2656 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2656 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2657 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2657 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2657 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2658 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2658 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2658 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2659 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2659 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2659 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2660 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2660 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2660 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2661 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2661 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2661 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2662 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2662 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2662 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2663 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2663 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2663 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2664 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2664 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2664 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2665 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2665 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2665 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2666 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2666 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2666 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2667 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2667 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2667 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2668 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2668 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2668 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2669 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2669 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2669 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2670 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2670 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2670 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2671 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2671 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2671 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2672 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2672 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2672 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2673 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2673 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2673 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2674 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2674 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2674 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2675 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2675 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2675 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2676 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2676 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2676 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2677 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2677 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2677 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2678 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2678 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2678 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2679 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2679 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2679 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2680 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2680 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2680 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2681 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2681 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2681 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2682 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2682 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2682 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2683 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2683 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2683 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2684 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2684 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2684 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2685 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2685 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2685 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2686 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2686 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2686 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2687 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2687 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2687 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2688 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2688 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2688 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2689 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2689 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2689 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2690 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2690 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2690 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2691 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2691 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2691 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2692 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2692 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2692 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2693 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2693 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2693 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2694 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2694 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2694 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2695 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2695 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2695 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2696 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2696 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2696 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2697 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2697 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2697 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2698 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2698 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2698 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2699 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2699 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2699 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2700 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2700 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2700 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2701 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2701 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2701 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2702 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2702 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2702 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2703 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2703 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2703 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2704 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2704 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2704 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2705 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2705 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2705 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2706 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2706 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2706 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2707 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2707 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2707 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2708 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2708 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2708 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2709 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2709 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2709 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2710 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2710 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2710 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2711 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2711 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2711 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2712 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2712 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2712 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2713 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2713 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2713 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2714 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2714 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2714 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2715 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2715 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2715 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2716 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2716 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2716 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2717 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2717 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2717 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2718 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2718 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2718 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2719 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'ha9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2719 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2719 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2720 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2720 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2720 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2721 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2721 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2721 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2722 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2722 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2722 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2723 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2723 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2723 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2724 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2724 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2724 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2725 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2725 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2725 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2726 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2726 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2726 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2727 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2727 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2727 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2728 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2728 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2728 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2729 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haa9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2729 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2729 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2730 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2730 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2730 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2731 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2731 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2731 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2732 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2732 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2732 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2733 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2733 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2733 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2734 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2734 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2734 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2735 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2735 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2735 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2736 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2736 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2736 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2737 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2737 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2737 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2738 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2738 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2738 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2739 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2739 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2739 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2740 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2740 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2740 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2741 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2741 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2741 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2742 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2742 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2742 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2743 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2743 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2743 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2744 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2744 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2744 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2745 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hab9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2745 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2745 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2746 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2746 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2746 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2747 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'habb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2747 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2747 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2748 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'habc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2748 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2748 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2749 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'habd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2749 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2749 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2750 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'habe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2750 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2750 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2751 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'habf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2751 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2751 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2752 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2752 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2752 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2753 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2753 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2753 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2754 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2754 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2754 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2755 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2755 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2755 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2756 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2756 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2756 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2757 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2757 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2757 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2758 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2758 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2758 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2759 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2759 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2759 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2760 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2760 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2760 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2761 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hac9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2761 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2761 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2762 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2762 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2762 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2763 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hacb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2763 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2763 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2764 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hacc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2764 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2764 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2765 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hacd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2765 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2765 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2766 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hace == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2766 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2766 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2767 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hacf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2767 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2767 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2768 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2768 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2768 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2769 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2769 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2769 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2770 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2770 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2770 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2771 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2771 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2771 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2772 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2772 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2772 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2773 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2773 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2773 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2774 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2774 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2774 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2775 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2775 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2775 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2776 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2776 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2776 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2777 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'had9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2777 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2777 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2778 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hada == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2778 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2778 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2779 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hadb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2779 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2779 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2780 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hadc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2780 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2780 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2781 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hadd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2781 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2781 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2782 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hade == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2782 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2782 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2783 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hadf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2783 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2783 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2784 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2784 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2784 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2785 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2785 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2785 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2786 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2786 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2786 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2787 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2787 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2787 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2788 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2788 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2788 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2789 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2789 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2789 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2790 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2790 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2790 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2791 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2791 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2791 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2792 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2792 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2792 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2793 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hae9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2793 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2793 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2794 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2794 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2794 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2795 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haeb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2795 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2795 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2796 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2796 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2796 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2797 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2797 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2797 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2798 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2798 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2798 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2799 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2799 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2799 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2800 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2800 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2800 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2801 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2801 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2801 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2802 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2802 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2802 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2803 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2803 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2803 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2804 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2804 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2804 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2805 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2805 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2805 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2806 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2806 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2806 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2807 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2807 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2807 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2808 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2808 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2808 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2809 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haf9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2809 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2809 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2810 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hafa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2810 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2810 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2811 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hafb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2811 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2811 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2812 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hafc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2812 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2812 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2813 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hafd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2813 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2813 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2814 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hafe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2814 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2814 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2815 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'haff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2815 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2815 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2816 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2816 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2816 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2817 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2817 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2817 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2818 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2818 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2818 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2819 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2819 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2819 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2820 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2820 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2820 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2821 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2821 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2821 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2822 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2822 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2822 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2823 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2823 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2823 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2824 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2824 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2824 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2825 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2825 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2825 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2826 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2826 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2826 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2827 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2827 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2827 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2828 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2828 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2828 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2829 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2829 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2829 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2830 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2830 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2830 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2831 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2831 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2831 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2832 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2832 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2832 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2833 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2833 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2833 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2834 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2834 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2834 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2835 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2835 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2835 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2836 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2836 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2836 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2837 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2837 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2837 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2838 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2838 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2838 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2839 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2839 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2839 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2840 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2840 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2840 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2841 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2841 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2841 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2842 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2842 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2842 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2843 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2843 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2843 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2844 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2844 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2844 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2845 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2845 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2845 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2846 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2846 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2846 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2847 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2847 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2847 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2848 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2848 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2848 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2849 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2849 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2849 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2850 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2850 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2850 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2851 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2851 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2851 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2852 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2852 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2852 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2853 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2853 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2853 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2854 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2854 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2854 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2855 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2855 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2855 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2856 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2856 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2856 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2857 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2857 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2857 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2858 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2858 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2858 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2859 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2859 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2859 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2860 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2860 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2860 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2861 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2861 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2861 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2862 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2862 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2862 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2863 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2863 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2863 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2864 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2864 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2864 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2865 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2865 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2865 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2866 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2866 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2866 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2867 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2867 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2867 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2868 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2868 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2868 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2869 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2869 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2869 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2870 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2870 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2870 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2871 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2871 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2871 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2872 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2872 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2872 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2873 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2873 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2873 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2874 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2874 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2874 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2875 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2875 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2875 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2876 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2876 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2876 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2877 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2877 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2877 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2878 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2878 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2878 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2879 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2879 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2879 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2880 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2880 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2880 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2881 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2881 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2881 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2882 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2882 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2882 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2883 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2883 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2883 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2884 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2884 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2884 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2885 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2885 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2885 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2886 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2886 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2886 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2887 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2887 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2887 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2888 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2888 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2888 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2889 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2889 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2889 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2890 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2890 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2890 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2891 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2891 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2891 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2892 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2892 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2892 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2893 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2893 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2893 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2894 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2894 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2894 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2895 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2895 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2895 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2896 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2896 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2896 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2897 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2897 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2897 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2898 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2898 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2898 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2899 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2899 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2899 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2900 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2900 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2900 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2901 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2901 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2901 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2902 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2902 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2902 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2903 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2903 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2903 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2904 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2904 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2904 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2905 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2905 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2905 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2906 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2906 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2906 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2907 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2907 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2907 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2908 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2908 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2908 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2909 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2909 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2909 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2910 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2910 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2910 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2911 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2911 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2911 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2912 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2912 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2912 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2913 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2913 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2913 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2914 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2914 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2914 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2915 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2915 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2915 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2916 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2916 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2916 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2917 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2917 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2917 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2918 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2918 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2918 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2919 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2919 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2919 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2920 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2920 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2920 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2921 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2921 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2921 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2922 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2922 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2922 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2923 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2923 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2923 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2924 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2924 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2924 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2925 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2925 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2925 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2926 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2926 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2926 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2927 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2927 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2927 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2928 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2928 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2928 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2929 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2929 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2929 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2930 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2930 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2930 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2931 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2931 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2931 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2932 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2932 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2932 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2933 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2933 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2933 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2934 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2934 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2934 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2935 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2935 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2935 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2936 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2936 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2936 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2937 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2937 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2937 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2938 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2938 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2938 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2939 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2939 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2939 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2940 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2940 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2940 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2941 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2941 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2941 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2942 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2942 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2942 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2943 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2943 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2943 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2944 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2944 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2944 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2945 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2945 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2945 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2946 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2946 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2946 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2947 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2947 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2947 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2948 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2948 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2948 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2949 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2949 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2949 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2950 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2950 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2950 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2951 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2951 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2951 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2952 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2952 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2952 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2953 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2953 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2953 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2954 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2954 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2954 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2955 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2955 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2955 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2956 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2956 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2956 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2957 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2957 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2957 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2958 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2958 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2958 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2959 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2959 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2959 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2960 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2960 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2960 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2961 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2961 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2961 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2962 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2962 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2962 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2963 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2963 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2963 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2964 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2964 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2964 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2965 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2965 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2965 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2966 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2966 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2966 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2967 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2967 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2967 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2968 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2968 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2968 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2969 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2969 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2969 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2970 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2970 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2970 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2971 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2971 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2971 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2972 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2972 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2972 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2973 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2973 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2973 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2974 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2974 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2974 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2975 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hb9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2975 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2975 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2976 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2976 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2976 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2977 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2977 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2977 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2978 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2978 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2978 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2979 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2979 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2979 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2980 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2980 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2980 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2981 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2981 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2981 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2982 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2982 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2982 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2983 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2983 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2983 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2984 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2984 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2984 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2985 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hba9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2985 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2985 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2986 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2986 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2986 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2987 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2987 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2987 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2988 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2988 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2988 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2989 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2989 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2989 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2990 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2990 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2990 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2991 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2991 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2991 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2992 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2992 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2992 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2993 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2993 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2993 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2994 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2994 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2994 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2995 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2995 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2995 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2996 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2996 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2996 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2997 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2997 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2997 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2998 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2998 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2998 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_2999 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_2999 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_2999 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3000 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3000 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3000 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3001 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3001 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3001 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3002 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3002 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3002 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3003 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbbb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3003 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3003 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3004 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbbc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3004 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3004 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3005 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbbd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3005 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3005 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3006 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbbe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3006 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3006 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3007 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbbf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3007 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3007 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3008 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3008 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3008 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3009 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3009 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3009 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3010 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3010 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3010 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3011 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3011 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3011 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3012 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3012 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3012 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3013 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3013 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3013 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3014 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3014 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3014 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3015 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3015 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3015 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3016 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3016 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3016 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3017 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbc9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3017 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3017 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3018 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3018 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3018 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3019 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbcb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3019 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3019 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3020 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbcc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3020 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3020 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3021 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbcd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3021 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3021 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3022 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3022 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3022 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3023 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbcf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3023 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3023 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3024 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3024 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3024 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3025 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3025 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3025 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3026 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3026 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3026 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3027 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3027 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3027 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3028 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3028 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3028 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3029 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3029 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3029 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3030 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3030 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3030 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3031 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3031 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3031 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3032 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3032 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3032 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3033 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbd9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3033 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3033 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3034 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3034 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3034 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3035 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbdb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3035 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3035 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3036 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbdc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3036 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3036 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3037 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbdd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3037 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3037 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3038 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbde == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3038 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3038 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3039 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbdf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3039 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3039 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3040 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3040 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3040 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3041 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3041 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3041 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3042 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3042 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3042 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3043 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3043 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3043 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3044 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3044 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3044 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3045 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3045 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3045 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3046 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3046 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3046 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3047 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3047 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3047 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3048 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3048 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3048 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3049 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbe9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3049 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3049 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3050 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3050 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3050 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3051 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbeb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3051 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3051 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3052 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3052 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3052 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3053 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3053 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3053 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3054 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3054 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3054 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3055 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3055 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3055 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3056 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3056 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3056 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3057 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3057 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3057 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3058 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3058 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3058 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3059 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3059 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3059 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3060 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3060 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3060 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3061 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3061 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3061 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3062 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3062 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3062 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3063 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3063 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3063 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3064 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3064 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3064 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3065 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbf9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3065 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3065 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3066 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbfa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3066 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3066 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3067 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbfb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3067 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3067 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3068 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbfc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3068 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3068 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3069 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbfd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3069 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3069 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3070 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbfe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3070 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3070 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3071 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hbff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3071 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3071 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3072 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3072 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3072 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3073 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3073 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3073 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3074 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3074 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3074 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3075 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3075 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3075 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3076 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3076 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3076 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3077 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3077 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3077 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3078 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3078 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3078 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3079 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3079 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3079 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3080 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3080 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3080 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3081 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3081 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3081 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3082 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3082 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3082 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3083 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3083 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3083 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3084 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3084 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3084 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3085 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3085 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3085 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3086 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3086 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3086 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3087 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3087 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3087 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3088 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3088 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3088 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3089 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3089 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3089 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3090 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3090 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3090 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3091 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3091 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3091 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3092 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3092 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3092 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3093 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3093 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3093 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3094 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3094 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3094 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3095 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3095 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3095 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3096 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3096 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3096 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3097 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3097 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3097 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3098 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3098 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3098 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3099 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3099 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3099 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3100 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3100 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3100 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3101 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3101 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3101 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3102 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3102 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3102 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3103 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3103 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3103 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3104 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3104 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3104 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3105 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3105 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3105 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3106 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3106 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3106 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3107 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3107 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3107 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3108 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3108 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3108 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3109 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3109 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3109 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3110 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3110 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3110 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3111 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3111 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3111 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3112 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3112 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3112 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3113 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3113 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3113 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3114 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3114 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3114 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3115 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3115 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3115 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3116 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3116 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3116 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3117 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3117 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3117 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3118 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3118 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3118 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3119 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3119 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3119 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3120 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3120 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3120 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3121 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3121 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3121 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3122 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3122 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3122 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3123 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3123 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3123 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3124 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3124 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3124 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3125 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3125 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3125 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3126 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3126 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3126 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3127 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3127 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3127 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3128 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3128 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3128 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3129 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3129 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3129 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3130 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3130 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3130 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3131 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3131 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3131 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3132 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3132 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3132 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3133 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3133 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3133 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3134 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3134 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3134 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3135 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3135 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3135 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3136 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3136 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3136 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3137 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3137 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3137 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3138 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3138 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3138 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3139 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3139 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3139 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3140 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3140 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3140 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3141 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3141 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3141 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3142 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3142 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3142 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3143 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3143 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3143 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3144 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3144 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3144 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3145 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3145 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3145 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3146 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3146 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3146 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3147 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3147 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3147 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3148 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3148 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3148 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3149 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3149 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3149 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3150 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3150 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3150 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3151 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3151 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3151 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3152 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3152 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3152 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3153 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3153 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3153 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3154 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3154 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3154 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3155 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3155 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3155 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3156 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3156 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3156 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3157 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3157 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3157 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3158 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3158 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3158 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3159 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3159 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3159 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3160 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3160 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3160 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3161 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3161 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3161 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3162 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3162 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3162 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3163 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3163 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3163 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3164 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3164 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3164 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3165 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3165 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3165 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3166 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3166 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3166 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3167 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3167 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3167 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3168 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3168 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3168 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3169 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3169 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3169 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3170 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3170 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3170 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3171 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3171 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3171 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3172 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3172 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3172 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3173 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3173 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3173 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3174 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3174 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3174 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3175 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3175 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3175 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3176 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3176 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3176 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3177 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3177 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3177 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3178 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3178 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3178 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3179 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3179 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3179 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3180 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3180 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3180 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3181 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3181 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3181 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3182 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3182 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3182 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3183 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3183 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3183 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3184 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3184 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3184 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3185 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3185 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3185 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3186 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3186 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3186 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3187 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3187 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3187 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3188 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3188 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3188 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3189 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3189 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3189 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3190 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3190 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3190 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3191 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3191 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3191 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3192 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3192 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3192 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3193 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3193 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3193 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3194 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3194 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3194 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3195 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3195 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3195 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3196 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3196 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3196 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3197 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3197 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3197 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3198 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3198 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3198 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3199 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3199 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3199 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3200 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3200 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3200 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3201 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3201 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3201 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3202 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3202 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3202 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3203 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3203 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3203 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3204 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3204 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3204 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3205 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3205 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3205 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3206 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3206 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3206 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3207 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3207 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3207 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3208 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3208 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3208 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3209 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3209 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3209 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3210 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3210 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3210 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3211 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3211 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3211 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3212 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3212 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3212 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3213 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3213 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3213 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3214 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3214 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3214 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3215 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3215 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3215 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3216 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3216 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3216 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3217 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3217 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3217 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3218 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3218 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3218 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3219 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3219 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3219 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3220 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3220 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3220 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3221 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3221 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3221 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3222 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3222 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3222 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3223 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3223 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3223 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3224 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3224 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3224 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3225 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3225 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3225 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3226 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3226 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3226 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3227 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3227 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3227 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3228 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3228 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3228 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3229 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3229 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3229 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3230 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3230 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3230 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3231 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hc9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3231 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3231 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3232 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3232 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3232 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3233 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3233 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3233 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3234 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3234 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3234 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3235 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3235 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3235 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3236 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3236 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3236 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3237 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3237 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3237 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3238 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3238 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3238 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3239 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3239 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3239 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3240 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3240 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3240 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3241 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hca9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3241 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3241 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3242 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3242 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3242 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3243 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3243 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3243 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3244 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3244 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3244 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3245 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3245 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3245 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3246 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3246 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3246 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3247 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3247 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3247 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3248 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3248 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3248 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3249 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3249 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3249 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3250 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3250 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3250 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3251 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3251 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3251 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3252 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3252 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3252 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3253 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3253 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3253 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3254 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3254 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3254 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3255 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3255 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3255 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3256 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3256 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3256 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3257 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3257 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3257 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3258 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3258 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3258 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3259 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcbb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3259 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3259 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3260 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcbc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3260 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3260 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3261 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcbd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3261 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3261 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3262 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcbe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3262 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3262 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3263 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcbf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3263 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3263 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3264 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3264 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3264 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3265 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3265 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3265 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3266 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3266 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3266 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3267 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3267 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3267 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3268 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3268 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3268 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3269 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3269 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3269 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3270 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3270 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3270 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3271 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3271 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3271 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3272 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3272 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3272 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3273 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcc9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3273 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3273 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3274 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3274 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3274 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3275 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hccb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3275 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3275 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3276 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hccc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3276 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3276 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3277 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hccd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3277 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3277 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3278 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3278 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3278 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3279 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hccf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3279 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3279 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3280 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3280 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3280 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3281 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3281 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3281 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3282 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3282 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3282 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3283 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3283 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3283 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3284 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3284 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3284 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3285 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3285 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3285 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3286 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3286 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3286 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3287 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3287 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3287 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3288 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3288 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3288 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3289 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcd9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3289 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3289 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3290 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3290 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3290 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3291 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcdb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3291 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3291 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3292 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcdc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3292 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3292 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3293 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcdd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3293 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3293 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3294 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcde == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3294 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3294 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3295 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcdf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3295 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3295 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3296 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3296 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3296 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3297 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3297 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3297 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3298 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3298 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3298 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3299 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3299 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3299 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3300 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3300 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3300 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3301 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3301 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3301 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3302 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3302 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3302 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3303 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3303 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3303 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3304 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3304 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3304 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3305 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hce9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3305 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3305 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3306 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3306 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3306 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3307 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hceb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3307 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3307 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3308 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3308 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3308 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3309 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hced == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3309 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3309 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3310 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3310 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3310 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3311 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3311 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3311 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3312 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3312 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3312 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3313 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3313 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3313 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3314 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3314 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3314 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3315 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3315 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3315 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3316 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3316 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3316 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3317 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3317 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3317 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3318 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3318 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3318 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3319 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3319 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3319 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3320 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3320 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3320 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3321 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcf9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3321 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3321 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3322 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcfa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3322 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3322 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3323 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcfb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3323 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3323 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3324 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcfc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3324 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3324 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3325 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcfd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3325 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3325 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3326 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcfe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3326 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3326 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3327 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hcff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3327 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3327 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3328 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3328 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3328 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3329 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3329 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3329 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3330 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3330 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3330 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3331 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3331 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3331 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3332 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3332 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3332 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3333 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3333 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3333 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3334 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3334 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3334 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3335 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3335 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3335 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3336 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3336 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3336 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3337 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3337 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3337 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3338 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3338 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3338 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3339 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3339 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3339 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3340 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3340 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3340 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3341 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3341 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3341 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3342 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3342 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3342 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3343 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3343 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3343 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3344 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3344 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3344 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3345 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3345 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3345 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3346 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3346 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3346 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3347 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3347 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3347 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3348 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3348 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3348 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3349 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3349 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3349 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3350 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3350 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3350 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3351 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3351 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3351 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3352 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3352 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3352 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3353 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3353 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3353 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3354 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3354 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3354 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3355 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3355 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3355 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3356 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3356 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3356 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3357 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3357 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3357 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3358 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3358 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3358 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3359 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3359 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3359 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3360 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3360 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3360 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3361 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3361 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3361 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3362 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3362 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3362 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3363 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3363 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3363 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3364 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3364 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3364 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3365 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3365 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3365 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3366 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3366 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3366 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3367 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3367 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3367 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3368 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3368 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3368 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3369 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3369 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3369 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3370 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3370 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3370 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3371 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3371 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3371 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3372 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3372 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3372 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3373 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3373 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3373 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3374 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3374 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3374 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3375 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3375 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3375 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3376 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3376 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3376 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3377 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3377 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3377 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3378 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3378 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3378 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3379 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3379 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3379 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3380 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3380 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3380 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3381 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3381 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3381 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3382 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3382 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3382 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3383 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3383 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3383 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3384 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3384 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3384 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3385 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3385 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3385 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3386 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3386 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3386 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3387 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3387 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3387 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3388 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3388 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3388 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3389 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3389 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3389 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3390 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3390 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3390 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3391 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3391 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3391 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3392 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3392 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3392 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3393 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3393 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3393 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3394 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3394 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3394 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3395 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3395 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3395 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3396 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3396 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3396 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3397 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3397 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3397 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3398 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3398 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3398 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3399 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3399 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3399 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3400 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3400 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3400 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3401 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3401 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3401 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3402 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3402 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3402 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3403 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3403 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3403 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3404 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3404 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3404 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3405 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3405 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3405 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3406 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3406 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3406 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3407 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3407 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3407 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3408 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3408 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3408 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3409 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3409 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3409 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3410 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3410 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3410 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3411 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3411 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3411 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3412 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3412 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3412 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3413 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3413 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3413 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3414 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3414 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3414 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3415 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3415 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3415 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3416 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3416 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3416 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3417 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3417 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3417 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3418 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3418 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3418 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3419 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3419 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3419 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3420 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3420 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3420 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3421 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3421 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3421 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3422 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3422 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3422 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3423 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3423 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3423 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3424 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3424 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3424 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3425 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3425 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3425 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3426 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3426 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3426 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3427 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3427 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3427 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3428 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3428 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3428 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3429 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3429 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3429 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3430 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3430 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3430 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3431 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3431 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3431 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3432 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3432 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3432 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3433 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3433 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3433 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3434 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3434 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3434 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3435 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3435 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3435 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3436 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3436 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3436 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3437 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3437 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3437 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3438 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3438 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3438 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3439 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3439 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3439 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3440 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3440 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3440 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3441 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3441 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3441 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3442 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3442 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3442 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3443 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3443 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3443 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3444 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3444 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3444 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3445 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3445 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3445 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3446 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3446 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3446 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3447 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3447 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3447 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3448 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3448 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3448 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3449 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3449 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3449 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3450 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3450 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3450 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3451 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3451 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3451 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3452 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3452 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3452 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3453 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3453 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3453 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3454 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3454 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3454 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3455 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3455 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3455 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3456 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3456 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3456 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3457 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3457 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3457 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3458 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3458 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3458 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3459 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3459 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3459 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3460 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3460 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3460 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3461 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3461 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3461 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3462 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3462 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3462 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3463 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3463 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3463 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3464 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3464 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3464 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3465 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3465 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3465 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3466 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3466 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3466 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3467 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3467 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3467 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3468 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3468 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3468 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3469 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3469 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3469 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3470 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3470 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3470 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3471 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3471 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3471 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3472 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3472 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3472 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3473 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3473 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3473 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3474 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3474 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3474 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3475 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3475 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3475 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3476 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3476 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3476 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3477 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3477 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3477 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3478 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3478 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3478 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3479 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3479 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3479 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3480 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3480 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3480 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3481 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3481 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3481 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3482 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3482 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3482 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3483 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3483 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3483 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3484 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3484 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3484 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3485 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3485 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3485 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3486 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3486 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3486 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3487 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hd9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3487 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3487 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3488 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3488 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3488 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3489 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3489 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3489 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3490 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3490 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3490 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3491 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3491 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3491 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3492 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3492 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3492 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3493 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3493 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3493 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3494 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3494 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3494 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3495 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3495 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3495 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3496 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3496 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3496 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3497 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hda9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3497 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3497 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3498 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3498 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3498 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3499 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3499 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3499 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3500 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3500 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3500 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3501 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3501 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3501 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3502 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3502 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3502 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3503 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3503 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3503 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3504 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3504 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3504 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3505 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3505 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3505 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3506 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3506 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3506 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3507 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3507 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3507 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3508 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3508 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3508 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3509 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3509 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3509 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3510 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3510 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3510 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3511 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3511 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3511 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3512 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3512 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3512 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3513 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3513 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3513 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3514 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3514 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3514 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3515 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdbb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3515 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3515 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3516 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdbc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3516 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3516 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3517 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdbd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3517 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3517 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3518 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdbe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3518 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3518 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3519 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdbf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3519 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3519 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3520 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3520 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3520 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3521 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3521 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3521 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3522 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3522 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3522 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3523 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3523 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3523 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3524 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3524 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3524 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3525 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3525 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3525 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3526 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3526 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3526 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3527 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3527 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3527 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3528 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3528 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3528 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3529 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdc9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3529 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3529 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3530 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3530 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3530 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3531 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdcb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3531 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3531 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3532 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdcc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3532 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3532 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3533 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdcd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3533 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3533 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3534 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3534 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3534 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3535 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdcf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3535 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3535 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3536 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3536 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3536 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3537 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3537 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3537 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3538 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3538 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3538 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3539 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3539 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3539 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3540 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3540 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3540 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3541 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3541 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3541 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3542 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3542 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3542 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3543 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3543 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3543 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3544 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3544 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3544 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3545 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdd9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3545 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3545 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3546 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3546 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3546 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3547 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hddb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3547 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3547 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3548 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hddc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3548 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3548 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3549 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hddd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3549 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3549 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3550 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdde == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3550 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3550 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3551 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hddf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3551 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3551 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3552 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3552 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3552 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3553 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3553 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3553 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3554 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3554 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3554 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3555 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3555 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3555 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3556 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3556 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3556 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3557 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3557 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3557 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3558 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3558 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3558 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3559 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3559 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3559 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3560 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3560 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3560 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3561 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hde9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3561 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3561 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3562 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3562 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3562 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3563 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdeb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3563 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3563 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3564 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3564 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3564 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3565 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hded == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3565 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3565 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3566 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3566 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3566 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3567 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3567 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3567 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3568 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3568 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3568 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3569 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3569 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3569 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3570 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3570 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3570 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3571 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3571 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3571 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3572 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3572 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3572 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3573 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3573 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3573 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3574 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3574 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3574 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3575 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3575 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3575 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3576 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3576 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3576 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3577 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdf9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3577 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3577 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3578 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdfa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3578 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3578 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3579 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdfb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3579 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3579 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3580 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdfc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3580 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3580 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3581 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdfd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3581 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3581 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3582 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdfe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3582 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3582 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3583 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hdff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3583 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3583 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3584 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3584 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3584 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3585 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3585 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3585 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3586 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3586 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3586 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3587 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3587 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3587 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3588 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3588 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3588 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3589 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3589 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3589 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3590 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3590 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3590 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3591 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3591 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3591 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3592 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3592 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3592 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3593 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3593 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3593 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3594 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3594 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3594 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3595 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3595 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3595 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3596 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3596 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3596 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3597 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3597 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3597 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3598 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3598 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3598 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3599 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3599 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3599 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3600 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3600 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3600 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3601 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3601 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3601 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3602 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3602 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3602 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3603 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3603 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3603 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3604 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3604 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3604 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3605 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3605 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3605 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3606 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3606 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3606 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3607 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3607 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3607 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3608 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3608 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3608 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3609 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3609 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3609 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3610 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3610 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3610 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3611 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3611 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3611 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3612 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3612 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3612 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3613 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3613 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3613 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3614 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3614 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3614 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3615 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3615 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3615 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3616 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3616 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3616 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3617 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3617 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3617 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3618 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3618 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3618 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3619 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3619 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3619 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3620 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3620 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3620 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3621 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3621 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3621 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3622 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3622 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3622 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3623 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3623 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3623 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3624 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3624 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3624 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3625 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3625 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3625 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3626 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3626 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3626 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3627 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3627 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3627 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3628 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3628 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3628 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3629 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3629 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3629 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3630 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3630 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3630 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3631 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3631 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3631 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3632 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3632 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3632 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3633 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3633 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3633 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3634 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3634 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3634 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3635 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3635 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3635 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3636 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3636 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3636 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3637 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3637 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3637 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3638 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3638 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3638 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3639 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3639 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3639 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3640 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3640 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3640 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3641 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3641 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3641 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3642 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3642 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3642 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3643 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3643 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3643 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3644 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3644 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3644 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3645 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3645 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3645 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3646 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3646 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3646 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3647 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3647 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3647 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3648 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3648 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3648 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3649 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3649 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3649 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3650 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3650 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3650 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3651 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3651 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3651 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3652 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3652 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3652 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3653 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3653 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3653 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3654 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3654 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3654 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3655 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3655 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3655 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3656 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3656 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3656 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3657 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3657 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3657 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3658 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3658 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3658 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3659 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3659 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3659 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3660 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3660 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3660 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3661 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3661 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3661 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3662 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3662 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3662 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3663 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3663 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3663 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3664 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3664 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3664 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3665 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3665 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3665 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3666 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3666 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3666 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3667 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3667 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3667 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3668 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3668 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3668 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3669 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3669 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3669 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3670 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3670 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3670 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3671 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3671 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3671 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3672 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3672 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3672 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3673 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3673 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3673 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3674 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3674 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3674 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3675 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3675 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3675 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3676 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3676 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3676 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3677 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3677 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3677 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3678 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3678 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3678 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3679 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3679 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3679 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3680 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3680 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3680 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3681 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3681 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3681 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3682 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3682 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3682 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3683 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3683 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3683 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3684 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3684 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3684 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3685 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3685 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3685 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3686 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3686 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3686 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3687 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3687 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3687 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3688 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3688 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3688 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3689 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3689 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3689 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3690 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3690 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3690 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3691 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3691 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3691 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3692 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3692 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3692 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3693 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3693 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3693 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3694 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3694 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3694 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3695 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3695 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3695 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3696 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3696 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3696 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3697 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3697 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3697 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3698 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3698 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3698 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3699 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3699 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3699 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3700 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3700 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3700 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3701 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3701 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3701 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3702 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3702 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3702 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3703 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3703 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3703 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3704 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3704 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3704 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3705 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3705 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3705 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3706 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3706 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3706 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3707 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3707 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3707 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3708 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3708 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3708 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3709 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3709 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3709 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3710 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3710 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3710 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3711 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3711 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3711 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3712 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3712 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3712 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3713 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3713 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3713 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3714 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3714 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3714 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3715 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3715 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3715 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3716 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3716 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3716 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3717 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3717 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3717 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3718 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3718 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3718 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3719 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3719 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3719 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3720 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3720 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3720 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3721 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3721 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3721 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3722 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3722 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3722 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3723 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3723 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3723 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3724 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3724 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3724 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3725 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3725 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3725 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3726 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3726 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3726 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3727 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3727 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3727 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3728 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3728 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3728 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3729 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3729 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3729 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3730 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3730 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3730 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3731 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3731 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3731 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3732 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3732 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3732 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3733 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3733 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3733 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3734 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3734 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3734 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3735 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3735 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3735 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3736 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3736 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3736 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3737 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3737 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3737 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3738 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3738 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3738 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3739 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3739 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3739 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3740 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3740 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3740 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3741 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3741 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3741 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3742 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3742 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3742 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3743 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'he9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3743 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3743 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3744 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3744 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3744 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3745 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3745 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3745 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3746 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3746 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3746 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3747 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3747 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3747 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3748 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3748 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3748 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3749 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3749 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3749 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3750 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3750 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3750 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3751 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3751 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3751 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3752 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3752 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3752 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3753 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hea9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3753 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3753 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3754 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3754 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3754 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3755 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3755 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3755 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3756 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3756 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3756 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3757 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'head == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3757 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3757 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3758 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3758 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3758 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3759 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3759 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3759 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3760 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3760 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3760 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3761 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3761 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3761 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3762 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3762 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3762 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3763 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3763 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3763 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3764 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3764 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3764 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3765 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3765 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3765 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3766 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3766 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3766 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3767 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3767 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3767 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3768 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3768 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3768 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3769 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3769 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3769 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3770 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3770 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3770 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3771 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hebb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3771 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3771 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3772 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hebc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3772 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3772 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3773 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hebd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3773 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3773 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3774 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hebe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3774 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3774 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3775 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hebf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3775 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3775 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3776 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3776 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3776 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3777 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3777 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3777 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3778 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3778 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3778 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3779 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3779 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3779 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3780 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3780 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3780 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3781 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3781 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3781 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3782 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3782 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3782 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3783 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3783 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3783 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3784 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3784 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3784 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3785 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hec9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3785 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3785 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3786 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3786 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3786 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3787 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hecb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3787 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3787 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3788 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hecc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3788 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3788 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3789 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hecd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3789 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3789 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3790 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hece == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3790 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3790 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3791 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hecf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3791 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3791 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3792 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3792 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3792 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3793 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3793 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3793 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3794 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3794 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3794 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3795 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3795 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3795 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3796 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3796 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3796 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3797 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3797 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3797 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3798 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3798 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3798 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3799 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3799 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3799 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3800 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3800 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3800 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3801 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hed9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3801 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3801 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3802 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3802 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3802 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3803 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hedb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3803 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3803 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3804 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hedc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3804 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3804 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3805 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hedd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3805 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3805 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3806 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hede == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3806 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3806 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3807 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hedf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3807 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3807 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3808 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3808 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3808 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3809 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3809 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3809 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3810 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3810 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3810 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3811 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3811 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3811 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3812 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3812 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3812 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3813 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3813 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3813 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3814 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3814 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3814 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3815 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3815 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3815 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3816 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3816 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3816 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3817 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hee9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3817 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3817 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3818 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3818 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3818 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3819 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heeb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3819 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3819 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3820 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3820 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3820 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3821 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3821 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3821 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3822 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3822 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3822 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3823 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3823 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3823 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3824 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3824 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3824 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3825 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3825 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3825 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3826 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3826 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3826 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3827 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3827 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3827 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3828 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3828 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3828 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3829 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3829 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3829 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3830 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3830 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3830 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3831 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3831 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3831 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3832 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3832 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3832 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3833 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hef9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3833 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3833 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3834 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hefa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3834 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3834 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3835 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hefb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3835 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3835 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3836 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hefc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3836 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3836 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3837 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hefd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3837 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3837 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3838 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hefe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3838 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3838 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3839 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'heff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3839 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3839 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3840 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf00 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3840 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3840 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3841 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf01 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3841 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3841 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3842 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf02 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3842 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3842 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3843 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf03 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3843 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3843 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3844 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf04 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3844 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3844 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3845 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf05 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3845 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3845 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3846 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf06 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3846 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3846 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3847 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf07 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3847 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3847 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3848 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf08 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3848 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3848 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3849 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf09 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3849 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3849 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3850 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3850 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3850 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3851 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3851 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3851 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3852 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3852 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3852 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3853 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3853 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3853 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3854 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3854 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3854 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3855 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf0f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3855 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3855 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3856 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf10 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3856 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3856 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3857 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf11 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3857 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3857 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3858 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf12 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3858 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3858 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3859 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf13 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3859 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3859 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3860 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf14 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3860 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3860 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3861 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf15 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3861 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3861 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3862 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf16 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3862 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3862 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3863 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf17 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3863 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3863 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3864 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf18 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3864 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3864 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3865 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf19 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3865 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3865 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3866 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3866 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3866 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3867 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3867 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3867 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3868 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3868 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3868 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3869 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3869 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3869 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3870 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3870 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3870 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3871 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf1f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3871 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3871 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3872 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf20 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3872 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3872 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3873 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf21 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3873 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3873 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3874 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf22 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3874 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3874 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3875 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf23 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3875 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3875 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3876 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf24 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3876 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3876 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3877 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf25 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3877 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3877 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3878 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf26 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3878 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3878 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3879 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf27 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3879 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3879 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3880 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf28 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3880 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3880 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3881 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf29 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3881 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3881 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3882 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3882 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3882 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3883 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3883 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3883 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3884 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3884 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3884 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3885 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3885 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3885 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3886 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3886 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3886 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3887 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf2f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3887 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3887 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3888 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf30 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3888 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3888 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3889 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf31 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3889 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3889 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3890 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf32 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3890 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3890 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3891 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf33 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3891 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3891 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3892 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf34 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3892 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3892 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3893 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf35 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3893 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3893 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3894 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf36 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3894 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3894 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3895 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf37 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3895 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3895 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3896 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf38 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3896 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3896 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3897 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf39 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3897 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3897 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3898 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3898 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3898 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3899 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3899 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3899 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3900 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3900 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3900 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3901 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3901 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3901 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3902 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3902 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3902 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3903 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf3f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3903 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3903 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3904 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf40 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3904 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3904 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3905 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf41 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3905 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3905 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3906 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf42 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3906 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3906 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3907 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf43 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3907 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3907 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3908 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf44 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3908 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3908 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3909 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf45 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3909 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3909 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3910 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf46 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3910 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3910 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3911 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf47 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3911 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3911 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3912 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf48 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3912 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3912 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3913 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf49 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3913 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3913 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3914 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3914 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3914 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3915 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3915 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3915 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3916 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3916 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3916 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3917 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3917 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3917 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3918 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3918 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3918 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3919 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf4f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3919 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3919 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3920 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf50 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3920 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3920 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3921 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf51 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3921 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3921 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3922 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf52 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3922 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3922 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3923 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf53 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3923 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3923 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3924 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf54 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3924 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3924 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3925 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf55 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3925 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3925 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3926 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf56 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3926 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3926 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3927 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf57 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3927 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3927 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3928 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf58 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3928 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3928 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3929 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf59 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3929 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3929 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3930 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3930 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3930 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3931 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3931 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3931 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3932 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3932 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3932 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3933 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3933 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3933 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3934 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3934 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3934 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3935 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf5f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3935 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3935 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3936 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf60 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3936 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3936 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3937 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf61 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3937 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3937 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3938 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf62 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3938 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3938 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3939 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf63 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3939 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3939 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3940 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf64 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3940 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3940 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3941 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf65 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3941 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3941 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3942 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf66 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3942 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3942 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3943 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf67 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3943 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3943 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3944 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf68 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3944 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3944 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3945 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf69 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3945 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3945 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3946 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3946 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3946 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3947 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3947 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3947 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3948 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3948 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3948 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3949 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3949 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3949 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3950 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3950 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3950 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3951 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf6f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3951 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3951 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3952 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf70 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3952 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3952 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3953 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf71 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3953 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3953 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3954 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf72 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3954 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3954 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3955 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf73 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3955 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3955 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3956 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf74 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3956 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3956 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3957 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf75 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3957 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3957 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3958 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf76 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3958 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3958 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3959 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf77 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3959 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3959 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3960 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf78 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3960 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3960 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3961 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf79 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3961 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3961 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3962 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3962 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3962 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3963 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3963 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3963 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3964 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3964 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3964 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3965 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3965 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3965 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3966 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3966 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3966 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3967 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf7f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3967 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3967 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3968 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf80 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3968 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3968 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3969 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf81 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3969 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3969 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3970 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf82 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3970 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3970 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3971 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf83 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3971 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3971 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3972 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf84 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3972 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3972 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3973 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf85 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3973 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3973 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3974 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf86 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3974 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3974 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3975 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf87 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3975 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3975 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3976 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf88 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3976 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3976 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3977 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf89 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3977 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3977 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3978 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3978 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3978 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3979 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3979 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3979 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3980 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3980 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3980 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3981 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3981 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3981 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3982 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3982 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3982 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3983 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf8f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3983 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3983 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3984 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf90 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3984 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3984 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3985 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf91 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3985 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3985 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3986 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf92 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3986 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3986 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3987 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf93 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3987 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3987 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3988 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf94 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3988 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3988 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3989 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf95 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3989 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3989 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3990 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf96 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3990 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3990 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3991 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf97 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3991 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3991 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3992 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf98 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3992 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3992 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3993 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf99 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3993 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3993 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3994 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9a == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3994 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3994 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3995 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9b == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3995 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3995 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3996 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9c == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3996 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3996 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3997 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9d == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3997 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3997 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3998 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9e == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3998 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3998 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_3999 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hf9f == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_3999 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_3999 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4000 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4000 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4000 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4001 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4001 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4001 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4002 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4002 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4002 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4003 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4003 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4003 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4004 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4004 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4004 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4005 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4005 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4005 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4006 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4006 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4006 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4007 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4007 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4007 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4008 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4008 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4008 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4009 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfa9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4009 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4009 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4010 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfaa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4010 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4010 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4011 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfab == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4011 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4011 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4012 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfac == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4012 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4012 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4013 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfad == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4013 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4013 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4014 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfae == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4014 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4014 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4015 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfaf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4015 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4015 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4016 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4016 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4016 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4017 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4017 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4017 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4018 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4018 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4018 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4019 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4019 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4019 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4020 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4020 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4020 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4021 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4021 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4021 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4022 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4022 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4022 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4023 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4023 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4023 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4024 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4024 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4024 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4025 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfb9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4025 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4025 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4026 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfba == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4026 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4026 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4027 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfbb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4027 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4027 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4028 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfbc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4028 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4028 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4029 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfbd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4029 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4029 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4030 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfbe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4030 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4030 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4031 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfbf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4031 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4031 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4032 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4032 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4032 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4033 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4033 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4033 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4034 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4034 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4034 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4035 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4035 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4035 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4036 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4036 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4036 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4037 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4037 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4037 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4038 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4038 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4038 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4039 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4039 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4039 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4040 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4040 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4040 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4041 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfc9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4041 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4041 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4042 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfca == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4042 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4042 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4043 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfcb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4043 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4043 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4044 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfcc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4044 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4044 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4045 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfcd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4045 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4045 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4046 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfce == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4046 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4046 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4047 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfcf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4047 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4047 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4048 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4048 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4048 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4049 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4049 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4049 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4050 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4050 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4050 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4051 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4051 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4051 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4052 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4052 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4052 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4053 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4053 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4053 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4054 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4054 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4054 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4055 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4055 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4055 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4056 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4056 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4056 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4057 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfd9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4057 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4057 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4058 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfda == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4058 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4058 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4059 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfdb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4059 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4059 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4060 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfdc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4060 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4060 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4061 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfdd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4061 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4061 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4062 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfde == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4062 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4062 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4063 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfdf == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4063 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4063 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4064 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4064 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4064 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4065 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4065 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4065 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4066 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4066 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4066 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4067 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4067 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4067 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4068 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4068 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4068 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4069 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4069 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4069 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4070 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4070 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4070 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4071 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4071 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4071 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4072 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4072 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4072 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4073 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfe9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4073 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4073 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4074 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfea == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4074 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4074 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4075 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfeb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4075 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4075 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4076 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfec == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4076 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4076 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4077 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfed == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4077 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4077 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4078 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfee == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4078 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4078 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4079 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfef == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4079 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4079 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4080 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff0 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4080 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4080 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4081 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff1 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4081 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4081 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4082 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff2 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4082 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4082 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4083 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff3 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4083 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4083 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4084 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff4 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4084 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4084 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4085 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff5 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4085 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4085 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4086 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff6 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4086 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4086 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4087 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff7 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4087 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4087 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4088 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff8 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4088 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4088 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4089 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hff9 == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4089 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4089 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4090 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hffa == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4090 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4090 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4091 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hffb == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4091 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4091 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4092 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hffc == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4092 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4092 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4093 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hffd == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4093 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4093 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4094 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hffe == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4094 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4094 <= _csr_wdata_T_9;
        end
      end
    end
    if (reset) begin // @[CSR.scala 31:26]
      reg_csr_4095 <= 32'h0; // @[CSR.scala 31:26]
    end else if (io_in_id_io_csr_cmd != 3'h0) begin // @[CSR.scala 49:31]
      if (12'hfff == csr_addr[11:0]) begin // @[CSR.scala 50:27]
        if (_csr_wdata_T) begin // @[Mux.scala 98:16]
          reg_csr_4095 <= io_in_id_io_op1_data;
        end else begin
          reg_csr_4095 <= _csr_wdata_T_9;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"csr_addr  = 0x%x\n",csr_addr); // @[CSR.scala 58:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"csr_rdata = 0x%x\n",_GEN_4095); // @[CSR.scala 59:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3) begin
          $fwrite(32'h80000002,"csr_wdata = 0x%x\n",csr_wdata); // @[CSR.scala 60:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_csr_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_csr_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_csr_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_csr_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_csr_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_csr_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_csr_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_csr_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_csr_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_csr_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_csr_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_csr_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_csr_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_csr_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_csr_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_csr_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_csr_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_csr_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_csr_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_csr_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_csr_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_csr_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_csr_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_csr_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_csr_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_csr_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_csr_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_csr_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_csr_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_csr_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_csr_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_csr_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  reg_csr_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  reg_csr_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  reg_csr_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  reg_csr_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_csr_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_csr_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_csr_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  reg_csr_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_csr_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  reg_csr_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  reg_csr_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  reg_csr_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  reg_csr_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  reg_csr_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  reg_csr_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  reg_csr_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_csr_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_csr_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  reg_csr_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  reg_csr_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  reg_csr_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  reg_csr_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  reg_csr_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  reg_csr_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  reg_csr_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  reg_csr_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  reg_csr_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  reg_csr_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  reg_csr_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  reg_csr_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  reg_csr_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  reg_csr_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  reg_csr_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  reg_csr_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  reg_csr_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  reg_csr_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  reg_csr_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  reg_csr_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  reg_csr_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  reg_csr_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  reg_csr_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  reg_csr_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  reg_csr_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  reg_csr_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  reg_csr_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  reg_csr_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  reg_csr_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  reg_csr_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  reg_csr_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  reg_csr_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  reg_csr_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  reg_csr_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  reg_csr_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  reg_csr_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  reg_csr_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  reg_csr_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  reg_csr_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  reg_csr_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  reg_csr_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  reg_csr_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  reg_csr_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  reg_csr_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  reg_csr_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  reg_csr_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  reg_csr_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  reg_csr_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  reg_csr_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  reg_csr_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  reg_csr_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  reg_csr_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  reg_csr_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  reg_csr_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  reg_csr_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  reg_csr_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  reg_csr_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  reg_csr_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  reg_csr_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  reg_csr_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  reg_csr_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  reg_csr_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  reg_csr_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  reg_csr_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  reg_csr_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  reg_csr_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  reg_csr_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  reg_csr_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  reg_csr_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  reg_csr_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  reg_csr_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  reg_csr_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  reg_csr_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  reg_csr_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  reg_csr_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  reg_csr_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  reg_csr_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  reg_csr_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  reg_csr_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  reg_csr_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  reg_csr_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  reg_csr_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  reg_csr_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  reg_csr_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  reg_csr_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  reg_csr_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  reg_csr_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  reg_csr_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  reg_csr_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  reg_csr_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  reg_csr_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  reg_csr_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  reg_csr_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  reg_csr_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  reg_csr_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  reg_csr_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  reg_csr_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  reg_csr_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  reg_csr_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  reg_csr_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  reg_csr_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  reg_csr_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  reg_csr_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  reg_csr_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  reg_csr_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  reg_csr_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  reg_csr_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  reg_csr_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  reg_csr_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  reg_csr_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  reg_csr_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  reg_csr_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  reg_csr_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  reg_csr_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  reg_csr_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  reg_csr_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  reg_csr_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  reg_csr_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  reg_csr_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  reg_csr_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  reg_csr_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  reg_csr_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  reg_csr_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  reg_csr_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  reg_csr_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  reg_csr_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  reg_csr_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  reg_csr_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  reg_csr_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  reg_csr_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  reg_csr_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  reg_csr_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  reg_csr_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  reg_csr_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  reg_csr_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  reg_csr_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  reg_csr_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  reg_csr_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  reg_csr_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  reg_csr_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  reg_csr_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  reg_csr_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  reg_csr_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  reg_csr_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  reg_csr_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  reg_csr_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  reg_csr_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  reg_csr_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  reg_csr_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  reg_csr_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  reg_csr_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  reg_csr_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  reg_csr_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  reg_csr_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  reg_csr_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  reg_csr_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  reg_csr_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  reg_csr_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  reg_csr_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  reg_csr_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  reg_csr_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  reg_csr_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  reg_csr_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  reg_csr_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  reg_csr_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  reg_csr_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  reg_csr_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  reg_csr_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  reg_csr_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  reg_csr_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  reg_csr_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  reg_csr_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  reg_csr_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  reg_csr_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  reg_csr_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  reg_csr_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  reg_csr_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  reg_csr_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  reg_csr_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  reg_csr_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  reg_csr_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  reg_csr_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  reg_csr_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  reg_csr_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  reg_csr_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  reg_csr_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  reg_csr_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  reg_csr_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  reg_csr_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  reg_csr_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  reg_csr_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  reg_csr_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  reg_csr_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  reg_csr_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  reg_csr_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  reg_csr_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  reg_csr_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  reg_csr_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  reg_csr_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  reg_csr_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  reg_csr_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  reg_csr_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  reg_csr_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  reg_csr_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  reg_csr_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  reg_csr_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  reg_csr_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  reg_csr_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  reg_csr_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  reg_csr_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  reg_csr_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  reg_csr_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  reg_csr_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  reg_csr_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  reg_csr_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  reg_csr_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  reg_csr_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  reg_csr_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  reg_csr_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  reg_csr_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  reg_csr_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  reg_csr_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  reg_csr_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  reg_csr_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  reg_csr_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  reg_csr_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  reg_csr_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  reg_csr_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  reg_csr_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  reg_csr_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  reg_csr_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  reg_csr_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  reg_csr_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  reg_csr_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  reg_csr_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  reg_csr_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  reg_csr_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  reg_csr_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  reg_csr_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  reg_csr_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  reg_csr_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  reg_csr_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  reg_csr_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  reg_csr_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  reg_csr_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  reg_csr_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  reg_csr_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  reg_csr_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  reg_csr_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  reg_csr_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  reg_csr_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  reg_csr_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  reg_csr_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  reg_csr_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  reg_csr_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  reg_csr_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  reg_csr_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  reg_csr_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  reg_csr_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  reg_csr_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  reg_csr_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  reg_csr_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  reg_csr_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  reg_csr_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  reg_csr_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  reg_csr_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  reg_csr_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  reg_csr_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  reg_csr_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  reg_csr_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  reg_csr_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  reg_csr_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  reg_csr_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  reg_csr_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  reg_csr_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  reg_csr_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  reg_csr_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  reg_csr_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  reg_csr_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  reg_csr_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  reg_csr_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  reg_csr_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  reg_csr_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  reg_csr_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  reg_csr_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  reg_csr_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  reg_csr_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  reg_csr_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  reg_csr_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  reg_csr_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  reg_csr_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  reg_csr_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  reg_csr_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  reg_csr_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  reg_csr_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  reg_csr_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  reg_csr_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  reg_csr_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  reg_csr_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  reg_csr_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  reg_csr_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  reg_csr_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  reg_csr_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  reg_csr_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  reg_csr_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  reg_csr_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  reg_csr_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  reg_csr_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  reg_csr_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  reg_csr_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  reg_csr_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  reg_csr_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  reg_csr_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  reg_csr_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  reg_csr_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  reg_csr_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  reg_csr_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  reg_csr_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  reg_csr_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  reg_csr_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  reg_csr_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  reg_csr_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  reg_csr_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  reg_csr_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  reg_csr_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  reg_csr_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  reg_csr_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  reg_csr_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  reg_csr_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  reg_csr_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  reg_csr_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  reg_csr_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  reg_csr_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  reg_csr_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  reg_csr_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  reg_csr_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  reg_csr_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  reg_csr_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  reg_csr_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  reg_csr_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  reg_csr_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  reg_csr_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  reg_csr_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  reg_csr_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  reg_csr_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  reg_csr_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  reg_csr_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  reg_csr_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  reg_csr_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  reg_csr_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  reg_csr_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  reg_csr_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  reg_csr_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  reg_csr_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  reg_csr_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  reg_csr_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  reg_csr_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  reg_csr_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  reg_csr_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  reg_csr_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  reg_csr_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  reg_csr_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  reg_csr_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  reg_csr_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  reg_csr_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  reg_csr_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  reg_csr_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  reg_csr_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  reg_csr_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  reg_csr_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  reg_csr_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  reg_csr_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  reg_csr_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  reg_csr_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  reg_csr_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  reg_csr_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  reg_csr_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  reg_csr_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  reg_csr_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  reg_csr_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  reg_csr_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  reg_csr_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  reg_csr_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  reg_csr_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  reg_csr_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  reg_csr_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  reg_csr_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  reg_csr_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  reg_csr_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  reg_csr_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  reg_csr_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  reg_csr_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  reg_csr_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  reg_csr_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  reg_csr_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  reg_csr_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  reg_csr_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  reg_csr_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  reg_csr_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  reg_csr_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  reg_csr_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  reg_csr_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  reg_csr_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  reg_csr_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  reg_csr_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  reg_csr_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  reg_csr_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  reg_csr_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  reg_csr_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  reg_csr_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  reg_csr_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  reg_csr_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  reg_csr_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  reg_csr_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  reg_csr_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  reg_csr_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  reg_csr_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  reg_csr_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  reg_csr_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  reg_csr_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  reg_csr_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  reg_csr_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  reg_csr_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  reg_csr_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  reg_csr_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  reg_csr_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  reg_csr_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  reg_csr_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  reg_csr_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  reg_csr_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  reg_csr_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  reg_csr_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  reg_csr_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  reg_csr_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  reg_csr_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  reg_csr_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  reg_csr_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  reg_csr_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  reg_csr_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  reg_csr_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  reg_csr_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  reg_csr_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  reg_csr_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  reg_csr_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  reg_csr_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  reg_csr_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  reg_csr_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  reg_csr_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  reg_csr_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  reg_csr_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  reg_csr_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  reg_csr_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  reg_csr_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  reg_csr_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  reg_csr_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  reg_csr_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  reg_csr_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  reg_csr_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  reg_csr_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  reg_csr_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  reg_csr_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  reg_csr_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  reg_csr_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  reg_csr_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  reg_csr_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  reg_csr_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  reg_csr_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  reg_csr_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  reg_csr_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  reg_csr_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  reg_csr_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  reg_csr_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  reg_csr_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  reg_csr_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  reg_csr_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  reg_csr_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  reg_csr_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  reg_csr_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  reg_csr_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  reg_csr_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  reg_csr_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  reg_csr_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  reg_csr_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  reg_csr_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  reg_csr_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  reg_csr_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  reg_csr_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  reg_csr_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  reg_csr_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  reg_csr_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  reg_csr_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  reg_csr_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  reg_csr_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  reg_csr_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  reg_csr_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  reg_csr_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  reg_csr_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  reg_csr_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  reg_csr_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  reg_csr_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  reg_csr_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  reg_csr_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  reg_csr_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  reg_csr_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  reg_csr_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  reg_csr_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  reg_csr_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  reg_csr_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  reg_csr_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  reg_csr_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  reg_csr_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  reg_csr_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  reg_csr_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  reg_csr_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  reg_csr_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  reg_csr_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  reg_csr_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  reg_csr_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  reg_csr_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  reg_csr_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  reg_csr_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  reg_csr_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  reg_csr_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  reg_csr_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  reg_csr_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  reg_csr_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  reg_csr_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  reg_csr_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  reg_csr_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  reg_csr_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  reg_csr_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  reg_csr_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  reg_csr_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  reg_csr_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  reg_csr_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  reg_csr_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  reg_csr_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  reg_csr_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  reg_csr_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  reg_csr_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  reg_csr_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  reg_csr_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  reg_csr_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  reg_csr_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  reg_csr_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  reg_csr_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  reg_csr_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  reg_csr_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  reg_csr_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  reg_csr_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  reg_csr_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  reg_csr_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  reg_csr_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  reg_csr_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  reg_csr_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  reg_csr_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  reg_csr_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  reg_csr_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  reg_csr_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  reg_csr_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  reg_csr_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  reg_csr_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  reg_csr_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  reg_csr_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  reg_csr_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  reg_csr_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  reg_csr_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  reg_csr_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  reg_csr_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  reg_csr_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  reg_csr_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  reg_csr_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  reg_csr_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  reg_csr_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  reg_csr_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  reg_csr_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  reg_csr_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  reg_csr_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  reg_csr_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  reg_csr_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  reg_csr_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  reg_csr_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  reg_csr_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  reg_csr_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  reg_csr_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  reg_csr_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  reg_csr_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  reg_csr_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  reg_csr_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  reg_csr_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  reg_csr_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  reg_csr_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  reg_csr_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  reg_csr_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  reg_csr_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  reg_csr_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  reg_csr_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  reg_csr_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  reg_csr_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  reg_csr_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  reg_csr_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  reg_csr_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  reg_csr_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  reg_csr_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  reg_csr_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  reg_csr_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  reg_csr_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  reg_csr_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  reg_csr_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  reg_csr_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  reg_csr_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  reg_csr_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  reg_csr_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  reg_csr_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  reg_csr_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  reg_csr_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  reg_csr_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  reg_csr_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  reg_csr_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  reg_csr_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  reg_csr_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  reg_csr_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  reg_csr_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  reg_csr_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  reg_csr_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  reg_csr_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  reg_csr_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  reg_csr_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  reg_csr_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  reg_csr_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  reg_csr_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  reg_csr_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  reg_csr_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  reg_csr_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  reg_csr_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  reg_csr_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  reg_csr_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  reg_csr_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  reg_csr_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  reg_csr_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  reg_csr_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  reg_csr_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  reg_csr_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  reg_csr_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  reg_csr_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  reg_csr_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  reg_csr_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  reg_csr_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  reg_csr_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  reg_csr_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  reg_csr_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  reg_csr_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  reg_csr_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  reg_csr_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  reg_csr_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  reg_csr_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  reg_csr_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  reg_csr_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  reg_csr_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  reg_csr_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  reg_csr_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  reg_csr_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  reg_csr_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  reg_csr_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  reg_csr_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  reg_csr_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  reg_csr_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  reg_csr_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  reg_csr_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  reg_csr_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  reg_csr_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  reg_csr_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  reg_csr_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  reg_csr_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  reg_csr_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  reg_csr_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  reg_csr_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  reg_csr_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  reg_csr_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  reg_csr_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  reg_csr_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  reg_csr_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  reg_csr_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  reg_csr_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  reg_csr_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  reg_csr_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  reg_csr_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  reg_csr_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  reg_csr_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  reg_csr_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  reg_csr_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  reg_csr_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  reg_csr_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  reg_csr_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  reg_csr_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  reg_csr_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  reg_csr_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  reg_csr_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  reg_csr_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  reg_csr_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  reg_csr_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  reg_csr_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  reg_csr_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  reg_csr_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  reg_csr_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  reg_csr_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  reg_csr_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  reg_csr_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  reg_csr_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  reg_csr_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  reg_csr_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  reg_csr_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  reg_csr_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  reg_csr_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  reg_csr_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  reg_csr_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  reg_csr_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  reg_csr_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  reg_csr_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  reg_csr_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  reg_csr_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  reg_csr_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  reg_csr_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  reg_csr_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  reg_csr_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  reg_csr_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  reg_csr_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  reg_csr_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  reg_csr_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  reg_csr_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  reg_csr_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  reg_csr_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  reg_csr_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  reg_csr_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  reg_csr_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  reg_csr_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  reg_csr_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  reg_csr_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  reg_csr_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  reg_csr_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  reg_csr_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  reg_csr_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  reg_csr_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  reg_csr_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  reg_csr_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  reg_csr_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  reg_csr_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  reg_csr_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  reg_csr_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  reg_csr_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  reg_csr_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  reg_csr_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  reg_csr_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  reg_csr_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  reg_csr_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  reg_csr_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  reg_csr_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  reg_csr_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  reg_csr_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  reg_csr_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  reg_csr_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  reg_csr_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  reg_csr_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  reg_csr_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  reg_csr_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  reg_csr_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  reg_csr_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  reg_csr_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  reg_csr_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  reg_csr_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  reg_csr_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  reg_csr_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  reg_csr_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  reg_csr_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  reg_csr_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  reg_csr_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  reg_csr_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  reg_csr_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  reg_csr_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  reg_csr_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  reg_csr_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  reg_csr_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  reg_csr_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  reg_csr_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  reg_csr_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  reg_csr_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  reg_csr_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  reg_csr_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  reg_csr_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  reg_csr_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  reg_csr_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  reg_csr_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  reg_csr_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  reg_csr_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  reg_csr_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  reg_csr_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  reg_csr_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  reg_csr_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  reg_csr_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  reg_csr_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  reg_csr_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  reg_csr_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  reg_csr_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  reg_csr_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  reg_csr_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  reg_csr_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  reg_csr_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  reg_csr_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  reg_csr_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  reg_csr_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  reg_csr_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  reg_csr_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  reg_csr_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  reg_csr_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  reg_csr_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  reg_csr_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  reg_csr_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  reg_csr_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  reg_csr_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  reg_csr_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  reg_csr_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  reg_csr_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  reg_csr_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  reg_csr_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  reg_csr_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  reg_csr_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  reg_csr_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  reg_csr_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  reg_csr_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  reg_csr_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  reg_csr_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  reg_csr_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  reg_csr_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  reg_csr_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  reg_csr_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  reg_csr_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  reg_csr_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  reg_csr_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  reg_csr_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  reg_csr_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  reg_csr_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  reg_csr_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  reg_csr_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  reg_csr_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  reg_csr_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  reg_csr_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  reg_csr_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  reg_csr_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  reg_csr_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  reg_csr_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  reg_csr_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  reg_csr_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  reg_csr_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  reg_csr_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  reg_csr_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  reg_csr_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  reg_csr_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  reg_csr_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  reg_csr_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  reg_csr_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  reg_csr_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  reg_csr_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  reg_csr_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  reg_csr_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  reg_csr_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  reg_csr_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  reg_csr_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  reg_csr_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  reg_csr_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  reg_csr_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  reg_csr_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  reg_csr_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  reg_csr_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  reg_csr_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  reg_csr_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  reg_csr_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  reg_csr_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  reg_csr_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  reg_csr_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  reg_csr_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  reg_csr_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  reg_csr_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  reg_csr_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  reg_csr_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  reg_csr_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  reg_csr_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  reg_csr_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  reg_csr_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  reg_csr_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  reg_csr_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  reg_csr_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  reg_csr_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  reg_csr_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  reg_csr_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  reg_csr_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  reg_csr_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  reg_csr_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  reg_csr_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  reg_csr_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  reg_csr_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  reg_csr_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  reg_csr_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  reg_csr_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  reg_csr_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  reg_csr_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  reg_csr_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  reg_csr_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  reg_csr_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  reg_csr_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  reg_csr_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  reg_csr_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  reg_csr_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  reg_csr_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  reg_csr_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  reg_csr_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  reg_csr_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  reg_csr_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  reg_csr_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  reg_csr_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  reg_csr_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  reg_csr_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  reg_csr_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  reg_csr_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  reg_csr_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  reg_csr_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  reg_csr_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  reg_csr_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  reg_csr_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  reg_csr_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  reg_csr_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  reg_csr_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  reg_csr_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  reg_csr_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  reg_csr_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  reg_csr_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  reg_csr_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  reg_csr_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  reg_csr_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  reg_csr_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  reg_csr_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  reg_csr_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  reg_csr_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  reg_csr_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  reg_csr_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  reg_csr_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  reg_csr_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  reg_csr_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  reg_csr_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  reg_csr_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  reg_csr_999 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  reg_csr_1000 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  reg_csr_1001 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  reg_csr_1002 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  reg_csr_1003 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  reg_csr_1004 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  reg_csr_1005 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  reg_csr_1006 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  reg_csr_1007 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  reg_csr_1008 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  reg_csr_1009 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  reg_csr_1010 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  reg_csr_1011 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  reg_csr_1012 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  reg_csr_1013 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  reg_csr_1014 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  reg_csr_1015 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  reg_csr_1016 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  reg_csr_1017 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  reg_csr_1018 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  reg_csr_1019 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  reg_csr_1020 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  reg_csr_1021 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  reg_csr_1022 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  reg_csr_1023 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  reg_csr_1024 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  reg_csr_1025 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  reg_csr_1026 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  reg_csr_1027 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  reg_csr_1028 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  reg_csr_1029 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  reg_csr_1030 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  reg_csr_1031 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  reg_csr_1032 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  reg_csr_1033 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  reg_csr_1034 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  reg_csr_1035 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  reg_csr_1036 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  reg_csr_1037 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  reg_csr_1038 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  reg_csr_1039 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  reg_csr_1040 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  reg_csr_1041 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  reg_csr_1042 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  reg_csr_1043 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  reg_csr_1044 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  reg_csr_1045 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  reg_csr_1046 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  reg_csr_1047 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  reg_csr_1048 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  reg_csr_1049 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  reg_csr_1050 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  reg_csr_1051 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  reg_csr_1052 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  reg_csr_1053 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  reg_csr_1054 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  reg_csr_1055 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  reg_csr_1056 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  reg_csr_1057 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  reg_csr_1058 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  reg_csr_1059 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  reg_csr_1060 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  reg_csr_1061 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  reg_csr_1062 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  reg_csr_1063 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  reg_csr_1064 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  reg_csr_1065 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  reg_csr_1066 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  reg_csr_1067 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  reg_csr_1068 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  reg_csr_1069 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  reg_csr_1070 = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  reg_csr_1071 = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  reg_csr_1072 = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  reg_csr_1073 = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  reg_csr_1074 = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  reg_csr_1075 = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  reg_csr_1076 = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  reg_csr_1077 = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  reg_csr_1078 = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  reg_csr_1079 = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  reg_csr_1080 = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  reg_csr_1081 = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  reg_csr_1082 = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  reg_csr_1083 = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  reg_csr_1084 = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  reg_csr_1085 = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  reg_csr_1086 = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  reg_csr_1087 = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  reg_csr_1088 = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  reg_csr_1089 = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  reg_csr_1090 = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  reg_csr_1091 = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  reg_csr_1092 = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  reg_csr_1093 = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  reg_csr_1094 = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  reg_csr_1095 = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  reg_csr_1096 = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  reg_csr_1097 = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  reg_csr_1098 = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  reg_csr_1099 = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  reg_csr_1100 = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  reg_csr_1101 = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  reg_csr_1102 = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  reg_csr_1103 = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  reg_csr_1104 = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  reg_csr_1105 = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  reg_csr_1106 = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  reg_csr_1107 = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  reg_csr_1108 = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  reg_csr_1109 = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  reg_csr_1110 = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  reg_csr_1111 = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  reg_csr_1112 = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  reg_csr_1113 = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  reg_csr_1114 = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  reg_csr_1115 = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  reg_csr_1116 = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  reg_csr_1117 = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  reg_csr_1118 = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  reg_csr_1119 = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  reg_csr_1120 = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  reg_csr_1121 = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  reg_csr_1122 = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  reg_csr_1123 = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  reg_csr_1124 = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  reg_csr_1125 = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  reg_csr_1126 = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  reg_csr_1127 = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  reg_csr_1128 = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  reg_csr_1129 = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  reg_csr_1130 = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  reg_csr_1131 = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  reg_csr_1132 = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  reg_csr_1133 = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  reg_csr_1134 = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  reg_csr_1135 = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  reg_csr_1136 = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  reg_csr_1137 = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  reg_csr_1138 = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  reg_csr_1139 = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  reg_csr_1140 = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  reg_csr_1141 = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  reg_csr_1142 = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  reg_csr_1143 = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  reg_csr_1144 = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  reg_csr_1145 = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  reg_csr_1146 = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  reg_csr_1147 = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  reg_csr_1148 = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  reg_csr_1149 = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  reg_csr_1150 = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  reg_csr_1151 = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  reg_csr_1152 = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  reg_csr_1153 = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  reg_csr_1154 = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  reg_csr_1155 = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  reg_csr_1156 = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  reg_csr_1157 = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  reg_csr_1158 = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  reg_csr_1159 = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  reg_csr_1160 = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  reg_csr_1161 = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  reg_csr_1162 = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  reg_csr_1163 = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  reg_csr_1164 = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  reg_csr_1165 = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  reg_csr_1166 = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  reg_csr_1167 = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  reg_csr_1168 = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  reg_csr_1169 = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  reg_csr_1170 = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  reg_csr_1171 = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  reg_csr_1172 = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  reg_csr_1173 = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  reg_csr_1174 = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  reg_csr_1175 = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  reg_csr_1176 = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  reg_csr_1177 = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  reg_csr_1178 = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  reg_csr_1179 = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  reg_csr_1180 = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  reg_csr_1181 = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  reg_csr_1182 = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  reg_csr_1183 = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  reg_csr_1184 = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  reg_csr_1185 = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  reg_csr_1186 = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  reg_csr_1187 = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  reg_csr_1188 = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  reg_csr_1189 = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  reg_csr_1190 = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  reg_csr_1191 = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  reg_csr_1192 = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  reg_csr_1193 = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  reg_csr_1194 = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  reg_csr_1195 = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  reg_csr_1196 = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  reg_csr_1197 = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  reg_csr_1198 = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  reg_csr_1199 = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  reg_csr_1200 = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  reg_csr_1201 = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  reg_csr_1202 = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  reg_csr_1203 = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  reg_csr_1204 = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  reg_csr_1205 = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  reg_csr_1206 = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  reg_csr_1207 = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  reg_csr_1208 = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  reg_csr_1209 = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  reg_csr_1210 = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  reg_csr_1211 = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  reg_csr_1212 = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  reg_csr_1213 = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  reg_csr_1214 = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  reg_csr_1215 = _RAND_1215[31:0];
  _RAND_1216 = {1{`RANDOM}};
  reg_csr_1216 = _RAND_1216[31:0];
  _RAND_1217 = {1{`RANDOM}};
  reg_csr_1217 = _RAND_1217[31:0];
  _RAND_1218 = {1{`RANDOM}};
  reg_csr_1218 = _RAND_1218[31:0];
  _RAND_1219 = {1{`RANDOM}};
  reg_csr_1219 = _RAND_1219[31:0];
  _RAND_1220 = {1{`RANDOM}};
  reg_csr_1220 = _RAND_1220[31:0];
  _RAND_1221 = {1{`RANDOM}};
  reg_csr_1221 = _RAND_1221[31:0];
  _RAND_1222 = {1{`RANDOM}};
  reg_csr_1222 = _RAND_1222[31:0];
  _RAND_1223 = {1{`RANDOM}};
  reg_csr_1223 = _RAND_1223[31:0];
  _RAND_1224 = {1{`RANDOM}};
  reg_csr_1224 = _RAND_1224[31:0];
  _RAND_1225 = {1{`RANDOM}};
  reg_csr_1225 = _RAND_1225[31:0];
  _RAND_1226 = {1{`RANDOM}};
  reg_csr_1226 = _RAND_1226[31:0];
  _RAND_1227 = {1{`RANDOM}};
  reg_csr_1227 = _RAND_1227[31:0];
  _RAND_1228 = {1{`RANDOM}};
  reg_csr_1228 = _RAND_1228[31:0];
  _RAND_1229 = {1{`RANDOM}};
  reg_csr_1229 = _RAND_1229[31:0];
  _RAND_1230 = {1{`RANDOM}};
  reg_csr_1230 = _RAND_1230[31:0];
  _RAND_1231 = {1{`RANDOM}};
  reg_csr_1231 = _RAND_1231[31:0];
  _RAND_1232 = {1{`RANDOM}};
  reg_csr_1232 = _RAND_1232[31:0];
  _RAND_1233 = {1{`RANDOM}};
  reg_csr_1233 = _RAND_1233[31:0];
  _RAND_1234 = {1{`RANDOM}};
  reg_csr_1234 = _RAND_1234[31:0];
  _RAND_1235 = {1{`RANDOM}};
  reg_csr_1235 = _RAND_1235[31:0];
  _RAND_1236 = {1{`RANDOM}};
  reg_csr_1236 = _RAND_1236[31:0];
  _RAND_1237 = {1{`RANDOM}};
  reg_csr_1237 = _RAND_1237[31:0];
  _RAND_1238 = {1{`RANDOM}};
  reg_csr_1238 = _RAND_1238[31:0];
  _RAND_1239 = {1{`RANDOM}};
  reg_csr_1239 = _RAND_1239[31:0];
  _RAND_1240 = {1{`RANDOM}};
  reg_csr_1240 = _RAND_1240[31:0];
  _RAND_1241 = {1{`RANDOM}};
  reg_csr_1241 = _RAND_1241[31:0];
  _RAND_1242 = {1{`RANDOM}};
  reg_csr_1242 = _RAND_1242[31:0];
  _RAND_1243 = {1{`RANDOM}};
  reg_csr_1243 = _RAND_1243[31:0];
  _RAND_1244 = {1{`RANDOM}};
  reg_csr_1244 = _RAND_1244[31:0];
  _RAND_1245 = {1{`RANDOM}};
  reg_csr_1245 = _RAND_1245[31:0];
  _RAND_1246 = {1{`RANDOM}};
  reg_csr_1246 = _RAND_1246[31:0];
  _RAND_1247 = {1{`RANDOM}};
  reg_csr_1247 = _RAND_1247[31:0];
  _RAND_1248 = {1{`RANDOM}};
  reg_csr_1248 = _RAND_1248[31:0];
  _RAND_1249 = {1{`RANDOM}};
  reg_csr_1249 = _RAND_1249[31:0];
  _RAND_1250 = {1{`RANDOM}};
  reg_csr_1250 = _RAND_1250[31:0];
  _RAND_1251 = {1{`RANDOM}};
  reg_csr_1251 = _RAND_1251[31:0];
  _RAND_1252 = {1{`RANDOM}};
  reg_csr_1252 = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  reg_csr_1253 = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  reg_csr_1254 = _RAND_1254[31:0];
  _RAND_1255 = {1{`RANDOM}};
  reg_csr_1255 = _RAND_1255[31:0];
  _RAND_1256 = {1{`RANDOM}};
  reg_csr_1256 = _RAND_1256[31:0];
  _RAND_1257 = {1{`RANDOM}};
  reg_csr_1257 = _RAND_1257[31:0];
  _RAND_1258 = {1{`RANDOM}};
  reg_csr_1258 = _RAND_1258[31:0];
  _RAND_1259 = {1{`RANDOM}};
  reg_csr_1259 = _RAND_1259[31:0];
  _RAND_1260 = {1{`RANDOM}};
  reg_csr_1260 = _RAND_1260[31:0];
  _RAND_1261 = {1{`RANDOM}};
  reg_csr_1261 = _RAND_1261[31:0];
  _RAND_1262 = {1{`RANDOM}};
  reg_csr_1262 = _RAND_1262[31:0];
  _RAND_1263 = {1{`RANDOM}};
  reg_csr_1263 = _RAND_1263[31:0];
  _RAND_1264 = {1{`RANDOM}};
  reg_csr_1264 = _RAND_1264[31:0];
  _RAND_1265 = {1{`RANDOM}};
  reg_csr_1265 = _RAND_1265[31:0];
  _RAND_1266 = {1{`RANDOM}};
  reg_csr_1266 = _RAND_1266[31:0];
  _RAND_1267 = {1{`RANDOM}};
  reg_csr_1267 = _RAND_1267[31:0];
  _RAND_1268 = {1{`RANDOM}};
  reg_csr_1268 = _RAND_1268[31:0];
  _RAND_1269 = {1{`RANDOM}};
  reg_csr_1269 = _RAND_1269[31:0];
  _RAND_1270 = {1{`RANDOM}};
  reg_csr_1270 = _RAND_1270[31:0];
  _RAND_1271 = {1{`RANDOM}};
  reg_csr_1271 = _RAND_1271[31:0];
  _RAND_1272 = {1{`RANDOM}};
  reg_csr_1272 = _RAND_1272[31:0];
  _RAND_1273 = {1{`RANDOM}};
  reg_csr_1273 = _RAND_1273[31:0];
  _RAND_1274 = {1{`RANDOM}};
  reg_csr_1274 = _RAND_1274[31:0];
  _RAND_1275 = {1{`RANDOM}};
  reg_csr_1275 = _RAND_1275[31:0];
  _RAND_1276 = {1{`RANDOM}};
  reg_csr_1276 = _RAND_1276[31:0];
  _RAND_1277 = {1{`RANDOM}};
  reg_csr_1277 = _RAND_1277[31:0];
  _RAND_1278 = {1{`RANDOM}};
  reg_csr_1278 = _RAND_1278[31:0];
  _RAND_1279 = {1{`RANDOM}};
  reg_csr_1279 = _RAND_1279[31:0];
  _RAND_1280 = {1{`RANDOM}};
  reg_csr_1280 = _RAND_1280[31:0];
  _RAND_1281 = {1{`RANDOM}};
  reg_csr_1281 = _RAND_1281[31:0];
  _RAND_1282 = {1{`RANDOM}};
  reg_csr_1282 = _RAND_1282[31:0];
  _RAND_1283 = {1{`RANDOM}};
  reg_csr_1283 = _RAND_1283[31:0];
  _RAND_1284 = {1{`RANDOM}};
  reg_csr_1284 = _RAND_1284[31:0];
  _RAND_1285 = {1{`RANDOM}};
  reg_csr_1285 = _RAND_1285[31:0];
  _RAND_1286 = {1{`RANDOM}};
  reg_csr_1286 = _RAND_1286[31:0];
  _RAND_1287 = {1{`RANDOM}};
  reg_csr_1287 = _RAND_1287[31:0];
  _RAND_1288 = {1{`RANDOM}};
  reg_csr_1288 = _RAND_1288[31:0];
  _RAND_1289 = {1{`RANDOM}};
  reg_csr_1289 = _RAND_1289[31:0];
  _RAND_1290 = {1{`RANDOM}};
  reg_csr_1290 = _RAND_1290[31:0];
  _RAND_1291 = {1{`RANDOM}};
  reg_csr_1291 = _RAND_1291[31:0];
  _RAND_1292 = {1{`RANDOM}};
  reg_csr_1292 = _RAND_1292[31:0];
  _RAND_1293 = {1{`RANDOM}};
  reg_csr_1293 = _RAND_1293[31:0];
  _RAND_1294 = {1{`RANDOM}};
  reg_csr_1294 = _RAND_1294[31:0];
  _RAND_1295 = {1{`RANDOM}};
  reg_csr_1295 = _RAND_1295[31:0];
  _RAND_1296 = {1{`RANDOM}};
  reg_csr_1296 = _RAND_1296[31:0];
  _RAND_1297 = {1{`RANDOM}};
  reg_csr_1297 = _RAND_1297[31:0];
  _RAND_1298 = {1{`RANDOM}};
  reg_csr_1298 = _RAND_1298[31:0];
  _RAND_1299 = {1{`RANDOM}};
  reg_csr_1299 = _RAND_1299[31:0];
  _RAND_1300 = {1{`RANDOM}};
  reg_csr_1300 = _RAND_1300[31:0];
  _RAND_1301 = {1{`RANDOM}};
  reg_csr_1301 = _RAND_1301[31:0];
  _RAND_1302 = {1{`RANDOM}};
  reg_csr_1302 = _RAND_1302[31:0];
  _RAND_1303 = {1{`RANDOM}};
  reg_csr_1303 = _RAND_1303[31:0];
  _RAND_1304 = {1{`RANDOM}};
  reg_csr_1304 = _RAND_1304[31:0];
  _RAND_1305 = {1{`RANDOM}};
  reg_csr_1305 = _RAND_1305[31:0];
  _RAND_1306 = {1{`RANDOM}};
  reg_csr_1306 = _RAND_1306[31:0];
  _RAND_1307 = {1{`RANDOM}};
  reg_csr_1307 = _RAND_1307[31:0];
  _RAND_1308 = {1{`RANDOM}};
  reg_csr_1308 = _RAND_1308[31:0];
  _RAND_1309 = {1{`RANDOM}};
  reg_csr_1309 = _RAND_1309[31:0];
  _RAND_1310 = {1{`RANDOM}};
  reg_csr_1310 = _RAND_1310[31:0];
  _RAND_1311 = {1{`RANDOM}};
  reg_csr_1311 = _RAND_1311[31:0];
  _RAND_1312 = {1{`RANDOM}};
  reg_csr_1312 = _RAND_1312[31:0];
  _RAND_1313 = {1{`RANDOM}};
  reg_csr_1313 = _RAND_1313[31:0];
  _RAND_1314 = {1{`RANDOM}};
  reg_csr_1314 = _RAND_1314[31:0];
  _RAND_1315 = {1{`RANDOM}};
  reg_csr_1315 = _RAND_1315[31:0];
  _RAND_1316 = {1{`RANDOM}};
  reg_csr_1316 = _RAND_1316[31:0];
  _RAND_1317 = {1{`RANDOM}};
  reg_csr_1317 = _RAND_1317[31:0];
  _RAND_1318 = {1{`RANDOM}};
  reg_csr_1318 = _RAND_1318[31:0];
  _RAND_1319 = {1{`RANDOM}};
  reg_csr_1319 = _RAND_1319[31:0];
  _RAND_1320 = {1{`RANDOM}};
  reg_csr_1320 = _RAND_1320[31:0];
  _RAND_1321 = {1{`RANDOM}};
  reg_csr_1321 = _RAND_1321[31:0];
  _RAND_1322 = {1{`RANDOM}};
  reg_csr_1322 = _RAND_1322[31:0];
  _RAND_1323 = {1{`RANDOM}};
  reg_csr_1323 = _RAND_1323[31:0];
  _RAND_1324 = {1{`RANDOM}};
  reg_csr_1324 = _RAND_1324[31:0];
  _RAND_1325 = {1{`RANDOM}};
  reg_csr_1325 = _RAND_1325[31:0];
  _RAND_1326 = {1{`RANDOM}};
  reg_csr_1326 = _RAND_1326[31:0];
  _RAND_1327 = {1{`RANDOM}};
  reg_csr_1327 = _RAND_1327[31:0];
  _RAND_1328 = {1{`RANDOM}};
  reg_csr_1328 = _RAND_1328[31:0];
  _RAND_1329 = {1{`RANDOM}};
  reg_csr_1329 = _RAND_1329[31:0];
  _RAND_1330 = {1{`RANDOM}};
  reg_csr_1330 = _RAND_1330[31:0];
  _RAND_1331 = {1{`RANDOM}};
  reg_csr_1331 = _RAND_1331[31:0];
  _RAND_1332 = {1{`RANDOM}};
  reg_csr_1332 = _RAND_1332[31:0];
  _RAND_1333 = {1{`RANDOM}};
  reg_csr_1333 = _RAND_1333[31:0];
  _RAND_1334 = {1{`RANDOM}};
  reg_csr_1334 = _RAND_1334[31:0];
  _RAND_1335 = {1{`RANDOM}};
  reg_csr_1335 = _RAND_1335[31:0];
  _RAND_1336 = {1{`RANDOM}};
  reg_csr_1336 = _RAND_1336[31:0];
  _RAND_1337 = {1{`RANDOM}};
  reg_csr_1337 = _RAND_1337[31:0];
  _RAND_1338 = {1{`RANDOM}};
  reg_csr_1338 = _RAND_1338[31:0];
  _RAND_1339 = {1{`RANDOM}};
  reg_csr_1339 = _RAND_1339[31:0];
  _RAND_1340 = {1{`RANDOM}};
  reg_csr_1340 = _RAND_1340[31:0];
  _RAND_1341 = {1{`RANDOM}};
  reg_csr_1341 = _RAND_1341[31:0];
  _RAND_1342 = {1{`RANDOM}};
  reg_csr_1342 = _RAND_1342[31:0];
  _RAND_1343 = {1{`RANDOM}};
  reg_csr_1343 = _RAND_1343[31:0];
  _RAND_1344 = {1{`RANDOM}};
  reg_csr_1344 = _RAND_1344[31:0];
  _RAND_1345 = {1{`RANDOM}};
  reg_csr_1345 = _RAND_1345[31:0];
  _RAND_1346 = {1{`RANDOM}};
  reg_csr_1346 = _RAND_1346[31:0];
  _RAND_1347 = {1{`RANDOM}};
  reg_csr_1347 = _RAND_1347[31:0];
  _RAND_1348 = {1{`RANDOM}};
  reg_csr_1348 = _RAND_1348[31:0];
  _RAND_1349 = {1{`RANDOM}};
  reg_csr_1349 = _RAND_1349[31:0];
  _RAND_1350 = {1{`RANDOM}};
  reg_csr_1350 = _RAND_1350[31:0];
  _RAND_1351 = {1{`RANDOM}};
  reg_csr_1351 = _RAND_1351[31:0];
  _RAND_1352 = {1{`RANDOM}};
  reg_csr_1352 = _RAND_1352[31:0];
  _RAND_1353 = {1{`RANDOM}};
  reg_csr_1353 = _RAND_1353[31:0];
  _RAND_1354 = {1{`RANDOM}};
  reg_csr_1354 = _RAND_1354[31:0];
  _RAND_1355 = {1{`RANDOM}};
  reg_csr_1355 = _RAND_1355[31:0];
  _RAND_1356 = {1{`RANDOM}};
  reg_csr_1356 = _RAND_1356[31:0];
  _RAND_1357 = {1{`RANDOM}};
  reg_csr_1357 = _RAND_1357[31:0];
  _RAND_1358 = {1{`RANDOM}};
  reg_csr_1358 = _RAND_1358[31:0];
  _RAND_1359 = {1{`RANDOM}};
  reg_csr_1359 = _RAND_1359[31:0];
  _RAND_1360 = {1{`RANDOM}};
  reg_csr_1360 = _RAND_1360[31:0];
  _RAND_1361 = {1{`RANDOM}};
  reg_csr_1361 = _RAND_1361[31:0];
  _RAND_1362 = {1{`RANDOM}};
  reg_csr_1362 = _RAND_1362[31:0];
  _RAND_1363 = {1{`RANDOM}};
  reg_csr_1363 = _RAND_1363[31:0];
  _RAND_1364 = {1{`RANDOM}};
  reg_csr_1364 = _RAND_1364[31:0];
  _RAND_1365 = {1{`RANDOM}};
  reg_csr_1365 = _RAND_1365[31:0];
  _RAND_1366 = {1{`RANDOM}};
  reg_csr_1366 = _RAND_1366[31:0];
  _RAND_1367 = {1{`RANDOM}};
  reg_csr_1367 = _RAND_1367[31:0];
  _RAND_1368 = {1{`RANDOM}};
  reg_csr_1368 = _RAND_1368[31:0];
  _RAND_1369 = {1{`RANDOM}};
  reg_csr_1369 = _RAND_1369[31:0];
  _RAND_1370 = {1{`RANDOM}};
  reg_csr_1370 = _RAND_1370[31:0];
  _RAND_1371 = {1{`RANDOM}};
  reg_csr_1371 = _RAND_1371[31:0];
  _RAND_1372 = {1{`RANDOM}};
  reg_csr_1372 = _RAND_1372[31:0];
  _RAND_1373 = {1{`RANDOM}};
  reg_csr_1373 = _RAND_1373[31:0];
  _RAND_1374 = {1{`RANDOM}};
  reg_csr_1374 = _RAND_1374[31:0];
  _RAND_1375 = {1{`RANDOM}};
  reg_csr_1375 = _RAND_1375[31:0];
  _RAND_1376 = {1{`RANDOM}};
  reg_csr_1376 = _RAND_1376[31:0];
  _RAND_1377 = {1{`RANDOM}};
  reg_csr_1377 = _RAND_1377[31:0];
  _RAND_1378 = {1{`RANDOM}};
  reg_csr_1378 = _RAND_1378[31:0];
  _RAND_1379 = {1{`RANDOM}};
  reg_csr_1379 = _RAND_1379[31:0];
  _RAND_1380 = {1{`RANDOM}};
  reg_csr_1380 = _RAND_1380[31:0];
  _RAND_1381 = {1{`RANDOM}};
  reg_csr_1381 = _RAND_1381[31:0];
  _RAND_1382 = {1{`RANDOM}};
  reg_csr_1382 = _RAND_1382[31:0];
  _RAND_1383 = {1{`RANDOM}};
  reg_csr_1383 = _RAND_1383[31:0];
  _RAND_1384 = {1{`RANDOM}};
  reg_csr_1384 = _RAND_1384[31:0];
  _RAND_1385 = {1{`RANDOM}};
  reg_csr_1385 = _RAND_1385[31:0];
  _RAND_1386 = {1{`RANDOM}};
  reg_csr_1386 = _RAND_1386[31:0];
  _RAND_1387 = {1{`RANDOM}};
  reg_csr_1387 = _RAND_1387[31:0];
  _RAND_1388 = {1{`RANDOM}};
  reg_csr_1388 = _RAND_1388[31:0];
  _RAND_1389 = {1{`RANDOM}};
  reg_csr_1389 = _RAND_1389[31:0];
  _RAND_1390 = {1{`RANDOM}};
  reg_csr_1390 = _RAND_1390[31:0];
  _RAND_1391 = {1{`RANDOM}};
  reg_csr_1391 = _RAND_1391[31:0];
  _RAND_1392 = {1{`RANDOM}};
  reg_csr_1392 = _RAND_1392[31:0];
  _RAND_1393 = {1{`RANDOM}};
  reg_csr_1393 = _RAND_1393[31:0];
  _RAND_1394 = {1{`RANDOM}};
  reg_csr_1394 = _RAND_1394[31:0];
  _RAND_1395 = {1{`RANDOM}};
  reg_csr_1395 = _RAND_1395[31:0];
  _RAND_1396 = {1{`RANDOM}};
  reg_csr_1396 = _RAND_1396[31:0];
  _RAND_1397 = {1{`RANDOM}};
  reg_csr_1397 = _RAND_1397[31:0];
  _RAND_1398 = {1{`RANDOM}};
  reg_csr_1398 = _RAND_1398[31:0];
  _RAND_1399 = {1{`RANDOM}};
  reg_csr_1399 = _RAND_1399[31:0];
  _RAND_1400 = {1{`RANDOM}};
  reg_csr_1400 = _RAND_1400[31:0];
  _RAND_1401 = {1{`RANDOM}};
  reg_csr_1401 = _RAND_1401[31:0];
  _RAND_1402 = {1{`RANDOM}};
  reg_csr_1402 = _RAND_1402[31:0];
  _RAND_1403 = {1{`RANDOM}};
  reg_csr_1403 = _RAND_1403[31:0];
  _RAND_1404 = {1{`RANDOM}};
  reg_csr_1404 = _RAND_1404[31:0];
  _RAND_1405 = {1{`RANDOM}};
  reg_csr_1405 = _RAND_1405[31:0];
  _RAND_1406 = {1{`RANDOM}};
  reg_csr_1406 = _RAND_1406[31:0];
  _RAND_1407 = {1{`RANDOM}};
  reg_csr_1407 = _RAND_1407[31:0];
  _RAND_1408 = {1{`RANDOM}};
  reg_csr_1408 = _RAND_1408[31:0];
  _RAND_1409 = {1{`RANDOM}};
  reg_csr_1409 = _RAND_1409[31:0];
  _RAND_1410 = {1{`RANDOM}};
  reg_csr_1410 = _RAND_1410[31:0];
  _RAND_1411 = {1{`RANDOM}};
  reg_csr_1411 = _RAND_1411[31:0];
  _RAND_1412 = {1{`RANDOM}};
  reg_csr_1412 = _RAND_1412[31:0];
  _RAND_1413 = {1{`RANDOM}};
  reg_csr_1413 = _RAND_1413[31:0];
  _RAND_1414 = {1{`RANDOM}};
  reg_csr_1414 = _RAND_1414[31:0];
  _RAND_1415 = {1{`RANDOM}};
  reg_csr_1415 = _RAND_1415[31:0];
  _RAND_1416 = {1{`RANDOM}};
  reg_csr_1416 = _RAND_1416[31:0];
  _RAND_1417 = {1{`RANDOM}};
  reg_csr_1417 = _RAND_1417[31:0];
  _RAND_1418 = {1{`RANDOM}};
  reg_csr_1418 = _RAND_1418[31:0];
  _RAND_1419 = {1{`RANDOM}};
  reg_csr_1419 = _RAND_1419[31:0];
  _RAND_1420 = {1{`RANDOM}};
  reg_csr_1420 = _RAND_1420[31:0];
  _RAND_1421 = {1{`RANDOM}};
  reg_csr_1421 = _RAND_1421[31:0];
  _RAND_1422 = {1{`RANDOM}};
  reg_csr_1422 = _RAND_1422[31:0];
  _RAND_1423 = {1{`RANDOM}};
  reg_csr_1423 = _RAND_1423[31:0];
  _RAND_1424 = {1{`RANDOM}};
  reg_csr_1424 = _RAND_1424[31:0];
  _RAND_1425 = {1{`RANDOM}};
  reg_csr_1425 = _RAND_1425[31:0];
  _RAND_1426 = {1{`RANDOM}};
  reg_csr_1426 = _RAND_1426[31:0];
  _RAND_1427 = {1{`RANDOM}};
  reg_csr_1427 = _RAND_1427[31:0];
  _RAND_1428 = {1{`RANDOM}};
  reg_csr_1428 = _RAND_1428[31:0];
  _RAND_1429 = {1{`RANDOM}};
  reg_csr_1429 = _RAND_1429[31:0];
  _RAND_1430 = {1{`RANDOM}};
  reg_csr_1430 = _RAND_1430[31:0];
  _RAND_1431 = {1{`RANDOM}};
  reg_csr_1431 = _RAND_1431[31:0];
  _RAND_1432 = {1{`RANDOM}};
  reg_csr_1432 = _RAND_1432[31:0];
  _RAND_1433 = {1{`RANDOM}};
  reg_csr_1433 = _RAND_1433[31:0];
  _RAND_1434 = {1{`RANDOM}};
  reg_csr_1434 = _RAND_1434[31:0];
  _RAND_1435 = {1{`RANDOM}};
  reg_csr_1435 = _RAND_1435[31:0];
  _RAND_1436 = {1{`RANDOM}};
  reg_csr_1436 = _RAND_1436[31:0];
  _RAND_1437 = {1{`RANDOM}};
  reg_csr_1437 = _RAND_1437[31:0];
  _RAND_1438 = {1{`RANDOM}};
  reg_csr_1438 = _RAND_1438[31:0];
  _RAND_1439 = {1{`RANDOM}};
  reg_csr_1439 = _RAND_1439[31:0];
  _RAND_1440 = {1{`RANDOM}};
  reg_csr_1440 = _RAND_1440[31:0];
  _RAND_1441 = {1{`RANDOM}};
  reg_csr_1441 = _RAND_1441[31:0];
  _RAND_1442 = {1{`RANDOM}};
  reg_csr_1442 = _RAND_1442[31:0];
  _RAND_1443 = {1{`RANDOM}};
  reg_csr_1443 = _RAND_1443[31:0];
  _RAND_1444 = {1{`RANDOM}};
  reg_csr_1444 = _RAND_1444[31:0];
  _RAND_1445 = {1{`RANDOM}};
  reg_csr_1445 = _RAND_1445[31:0];
  _RAND_1446 = {1{`RANDOM}};
  reg_csr_1446 = _RAND_1446[31:0];
  _RAND_1447 = {1{`RANDOM}};
  reg_csr_1447 = _RAND_1447[31:0];
  _RAND_1448 = {1{`RANDOM}};
  reg_csr_1448 = _RAND_1448[31:0];
  _RAND_1449 = {1{`RANDOM}};
  reg_csr_1449 = _RAND_1449[31:0];
  _RAND_1450 = {1{`RANDOM}};
  reg_csr_1450 = _RAND_1450[31:0];
  _RAND_1451 = {1{`RANDOM}};
  reg_csr_1451 = _RAND_1451[31:0];
  _RAND_1452 = {1{`RANDOM}};
  reg_csr_1452 = _RAND_1452[31:0];
  _RAND_1453 = {1{`RANDOM}};
  reg_csr_1453 = _RAND_1453[31:0];
  _RAND_1454 = {1{`RANDOM}};
  reg_csr_1454 = _RAND_1454[31:0];
  _RAND_1455 = {1{`RANDOM}};
  reg_csr_1455 = _RAND_1455[31:0];
  _RAND_1456 = {1{`RANDOM}};
  reg_csr_1456 = _RAND_1456[31:0];
  _RAND_1457 = {1{`RANDOM}};
  reg_csr_1457 = _RAND_1457[31:0];
  _RAND_1458 = {1{`RANDOM}};
  reg_csr_1458 = _RAND_1458[31:0];
  _RAND_1459 = {1{`RANDOM}};
  reg_csr_1459 = _RAND_1459[31:0];
  _RAND_1460 = {1{`RANDOM}};
  reg_csr_1460 = _RAND_1460[31:0];
  _RAND_1461 = {1{`RANDOM}};
  reg_csr_1461 = _RAND_1461[31:0];
  _RAND_1462 = {1{`RANDOM}};
  reg_csr_1462 = _RAND_1462[31:0];
  _RAND_1463 = {1{`RANDOM}};
  reg_csr_1463 = _RAND_1463[31:0];
  _RAND_1464 = {1{`RANDOM}};
  reg_csr_1464 = _RAND_1464[31:0];
  _RAND_1465 = {1{`RANDOM}};
  reg_csr_1465 = _RAND_1465[31:0];
  _RAND_1466 = {1{`RANDOM}};
  reg_csr_1466 = _RAND_1466[31:0];
  _RAND_1467 = {1{`RANDOM}};
  reg_csr_1467 = _RAND_1467[31:0];
  _RAND_1468 = {1{`RANDOM}};
  reg_csr_1468 = _RAND_1468[31:0];
  _RAND_1469 = {1{`RANDOM}};
  reg_csr_1469 = _RAND_1469[31:0];
  _RAND_1470 = {1{`RANDOM}};
  reg_csr_1470 = _RAND_1470[31:0];
  _RAND_1471 = {1{`RANDOM}};
  reg_csr_1471 = _RAND_1471[31:0];
  _RAND_1472 = {1{`RANDOM}};
  reg_csr_1472 = _RAND_1472[31:0];
  _RAND_1473 = {1{`RANDOM}};
  reg_csr_1473 = _RAND_1473[31:0];
  _RAND_1474 = {1{`RANDOM}};
  reg_csr_1474 = _RAND_1474[31:0];
  _RAND_1475 = {1{`RANDOM}};
  reg_csr_1475 = _RAND_1475[31:0];
  _RAND_1476 = {1{`RANDOM}};
  reg_csr_1476 = _RAND_1476[31:0];
  _RAND_1477 = {1{`RANDOM}};
  reg_csr_1477 = _RAND_1477[31:0];
  _RAND_1478 = {1{`RANDOM}};
  reg_csr_1478 = _RAND_1478[31:0];
  _RAND_1479 = {1{`RANDOM}};
  reg_csr_1479 = _RAND_1479[31:0];
  _RAND_1480 = {1{`RANDOM}};
  reg_csr_1480 = _RAND_1480[31:0];
  _RAND_1481 = {1{`RANDOM}};
  reg_csr_1481 = _RAND_1481[31:0];
  _RAND_1482 = {1{`RANDOM}};
  reg_csr_1482 = _RAND_1482[31:0];
  _RAND_1483 = {1{`RANDOM}};
  reg_csr_1483 = _RAND_1483[31:0];
  _RAND_1484 = {1{`RANDOM}};
  reg_csr_1484 = _RAND_1484[31:0];
  _RAND_1485 = {1{`RANDOM}};
  reg_csr_1485 = _RAND_1485[31:0];
  _RAND_1486 = {1{`RANDOM}};
  reg_csr_1486 = _RAND_1486[31:0];
  _RAND_1487 = {1{`RANDOM}};
  reg_csr_1487 = _RAND_1487[31:0];
  _RAND_1488 = {1{`RANDOM}};
  reg_csr_1488 = _RAND_1488[31:0];
  _RAND_1489 = {1{`RANDOM}};
  reg_csr_1489 = _RAND_1489[31:0];
  _RAND_1490 = {1{`RANDOM}};
  reg_csr_1490 = _RAND_1490[31:0];
  _RAND_1491 = {1{`RANDOM}};
  reg_csr_1491 = _RAND_1491[31:0];
  _RAND_1492 = {1{`RANDOM}};
  reg_csr_1492 = _RAND_1492[31:0];
  _RAND_1493 = {1{`RANDOM}};
  reg_csr_1493 = _RAND_1493[31:0];
  _RAND_1494 = {1{`RANDOM}};
  reg_csr_1494 = _RAND_1494[31:0];
  _RAND_1495 = {1{`RANDOM}};
  reg_csr_1495 = _RAND_1495[31:0];
  _RAND_1496 = {1{`RANDOM}};
  reg_csr_1496 = _RAND_1496[31:0];
  _RAND_1497 = {1{`RANDOM}};
  reg_csr_1497 = _RAND_1497[31:0];
  _RAND_1498 = {1{`RANDOM}};
  reg_csr_1498 = _RAND_1498[31:0];
  _RAND_1499 = {1{`RANDOM}};
  reg_csr_1499 = _RAND_1499[31:0];
  _RAND_1500 = {1{`RANDOM}};
  reg_csr_1500 = _RAND_1500[31:0];
  _RAND_1501 = {1{`RANDOM}};
  reg_csr_1501 = _RAND_1501[31:0];
  _RAND_1502 = {1{`RANDOM}};
  reg_csr_1502 = _RAND_1502[31:0];
  _RAND_1503 = {1{`RANDOM}};
  reg_csr_1503 = _RAND_1503[31:0];
  _RAND_1504 = {1{`RANDOM}};
  reg_csr_1504 = _RAND_1504[31:0];
  _RAND_1505 = {1{`RANDOM}};
  reg_csr_1505 = _RAND_1505[31:0];
  _RAND_1506 = {1{`RANDOM}};
  reg_csr_1506 = _RAND_1506[31:0];
  _RAND_1507 = {1{`RANDOM}};
  reg_csr_1507 = _RAND_1507[31:0];
  _RAND_1508 = {1{`RANDOM}};
  reg_csr_1508 = _RAND_1508[31:0];
  _RAND_1509 = {1{`RANDOM}};
  reg_csr_1509 = _RAND_1509[31:0];
  _RAND_1510 = {1{`RANDOM}};
  reg_csr_1510 = _RAND_1510[31:0];
  _RAND_1511 = {1{`RANDOM}};
  reg_csr_1511 = _RAND_1511[31:0];
  _RAND_1512 = {1{`RANDOM}};
  reg_csr_1512 = _RAND_1512[31:0];
  _RAND_1513 = {1{`RANDOM}};
  reg_csr_1513 = _RAND_1513[31:0];
  _RAND_1514 = {1{`RANDOM}};
  reg_csr_1514 = _RAND_1514[31:0];
  _RAND_1515 = {1{`RANDOM}};
  reg_csr_1515 = _RAND_1515[31:0];
  _RAND_1516 = {1{`RANDOM}};
  reg_csr_1516 = _RAND_1516[31:0];
  _RAND_1517 = {1{`RANDOM}};
  reg_csr_1517 = _RAND_1517[31:0];
  _RAND_1518 = {1{`RANDOM}};
  reg_csr_1518 = _RAND_1518[31:0];
  _RAND_1519 = {1{`RANDOM}};
  reg_csr_1519 = _RAND_1519[31:0];
  _RAND_1520 = {1{`RANDOM}};
  reg_csr_1520 = _RAND_1520[31:0];
  _RAND_1521 = {1{`RANDOM}};
  reg_csr_1521 = _RAND_1521[31:0];
  _RAND_1522 = {1{`RANDOM}};
  reg_csr_1522 = _RAND_1522[31:0];
  _RAND_1523 = {1{`RANDOM}};
  reg_csr_1523 = _RAND_1523[31:0];
  _RAND_1524 = {1{`RANDOM}};
  reg_csr_1524 = _RAND_1524[31:0];
  _RAND_1525 = {1{`RANDOM}};
  reg_csr_1525 = _RAND_1525[31:0];
  _RAND_1526 = {1{`RANDOM}};
  reg_csr_1526 = _RAND_1526[31:0];
  _RAND_1527 = {1{`RANDOM}};
  reg_csr_1527 = _RAND_1527[31:0];
  _RAND_1528 = {1{`RANDOM}};
  reg_csr_1528 = _RAND_1528[31:0];
  _RAND_1529 = {1{`RANDOM}};
  reg_csr_1529 = _RAND_1529[31:0];
  _RAND_1530 = {1{`RANDOM}};
  reg_csr_1530 = _RAND_1530[31:0];
  _RAND_1531 = {1{`RANDOM}};
  reg_csr_1531 = _RAND_1531[31:0];
  _RAND_1532 = {1{`RANDOM}};
  reg_csr_1532 = _RAND_1532[31:0];
  _RAND_1533 = {1{`RANDOM}};
  reg_csr_1533 = _RAND_1533[31:0];
  _RAND_1534 = {1{`RANDOM}};
  reg_csr_1534 = _RAND_1534[31:0];
  _RAND_1535 = {1{`RANDOM}};
  reg_csr_1535 = _RAND_1535[31:0];
  _RAND_1536 = {1{`RANDOM}};
  reg_csr_1536 = _RAND_1536[31:0];
  _RAND_1537 = {1{`RANDOM}};
  reg_csr_1537 = _RAND_1537[31:0];
  _RAND_1538 = {1{`RANDOM}};
  reg_csr_1538 = _RAND_1538[31:0];
  _RAND_1539 = {1{`RANDOM}};
  reg_csr_1539 = _RAND_1539[31:0];
  _RAND_1540 = {1{`RANDOM}};
  reg_csr_1540 = _RAND_1540[31:0];
  _RAND_1541 = {1{`RANDOM}};
  reg_csr_1541 = _RAND_1541[31:0];
  _RAND_1542 = {1{`RANDOM}};
  reg_csr_1542 = _RAND_1542[31:0];
  _RAND_1543 = {1{`RANDOM}};
  reg_csr_1543 = _RAND_1543[31:0];
  _RAND_1544 = {1{`RANDOM}};
  reg_csr_1544 = _RAND_1544[31:0];
  _RAND_1545 = {1{`RANDOM}};
  reg_csr_1545 = _RAND_1545[31:0];
  _RAND_1546 = {1{`RANDOM}};
  reg_csr_1546 = _RAND_1546[31:0];
  _RAND_1547 = {1{`RANDOM}};
  reg_csr_1547 = _RAND_1547[31:0];
  _RAND_1548 = {1{`RANDOM}};
  reg_csr_1548 = _RAND_1548[31:0];
  _RAND_1549 = {1{`RANDOM}};
  reg_csr_1549 = _RAND_1549[31:0];
  _RAND_1550 = {1{`RANDOM}};
  reg_csr_1550 = _RAND_1550[31:0];
  _RAND_1551 = {1{`RANDOM}};
  reg_csr_1551 = _RAND_1551[31:0];
  _RAND_1552 = {1{`RANDOM}};
  reg_csr_1552 = _RAND_1552[31:0];
  _RAND_1553 = {1{`RANDOM}};
  reg_csr_1553 = _RAND_1553[31:0];
  _RAND_1554 = {1{`RANDOM}};
  reg_csr_1554 = _RAND_1554[31:0];
  _RAND_1555 = {1{`RANDOM}};
  reg_csr_1555 = _RAND_1555[31:0];
  _RAND_1556 = {1{`RANDOM}};
  reg_csr_1556 = _RAND_1556[31:0];
  _RAND_1557 = {1{`RANDOM}};
  reg_csr_1557 = _RAND_1557[31:0];
  _RAND_1558 = {1{`RANDOM}};
  reg_csr_1558 = _RAND_1558[31:0];
  _RAND_1559 = {1{`RANDOM}};
  reg_csr_1559 = _RAND_1559[31:0];
  _RAND_1560 = {1{`RANDOM}};
  reg_csr_1560 = _RAND_1560[31:0];
  _RAND_1561 = {1{`RANDOM}};
  reg_csr_1561 = _RAND_1561[31:0];
  _RAND_1562 = {1{`RANDOM}};
  reg_csr_1562 = _RAND_1562[31:0];
  _RAND_1563 = {1{`RANDOM}};
  reg_csr_1563 = _RAND_1563[31:0];
  _RAND_1564 = {1{`RANDOM}};
  reg_csr_1564 = _RAND_1564[31:0];
  _RAND_1565 = {1{`RANDOM}};
  reg_csr_1565 = _RAND_1565[31:0];
  _RAND_1566 = {1{`RANDOM}};
  reg_csr_1566 = _RAND_1566[31:0];
  _RAND_1567 = {1{`RANDOM}};
  reg_csr_1567 = _RAND_1567[31:0];
  _RAND_1568 = {1{`RANDOM}};
  reg_csr_1568 = _RAND_1568[31:0];
  _RAND_1569 = {1{`RANDOM}};
  reg_csr_1569 = _RAND_1569[31:0];
  _RAND_1570 = {1{`RANDOM}};
  reg_csr_1570 = _RAND_1570[31:0];
  _RAND_1571 = {1{`RANDOM}};
  reg_csr_1571 = _RAND_1571[31:0];
  _RAND_1572 = {1{`RANDOM}};
  reg_csr_1572 = _RAND_1572[31:0];
  _RAND_1573 = {1{`RANDOM}};
  reg_csr_1573 = _RAND_1573[31:0];
  _RAND_1574 = {1{`RANDOM}};
  reg_csr_1574 = _RAND_1574[31:0];
  _RAND_1575 = {1{`RANDOM}};
  reg_csr_1575 = _RAND_1575[31:0];
  _RAND_1576 = {1{`RANDOM}};
  reg_csr_1576 = _RAND_1576[31:0];
  _RAND_1577 = {1{`RANDOM}};
  reg_csr_1577 = _RAND_1577[31:0];
  _RAND_1578 = {1{`RANDOM}};
  reg_csr_1578 = _RAND_1578[31:0];
  _RAND_1579 = {1{`RANDOM}};
  reg_csr_1579 = _RAND_1579[31:0];
  _RAND_1580 = {1{`RANDOM}};
  reg_csr_1580 = _RAND_1580[31:0];
  _RAND_1581 = {1{`RANDOM}};
  reg_csr_1581 = _RAND_1581[31:0];
  _RAND_1582 = {1{`RANDOM}};
  reg_csr_1582 = _RAND_1582[31:0];
  _RAND_1583 = {1{`RANDOM}};
  reg_csr_1583 = _RAND_1583[31:0];
  _RAND_1584 = {1{`RANDOM}};
  reg_csr_1584 = _RAND_1584[31:0];
  _RAND_1585 = {1{`RANDOM}};
  reg_csr_1585 = _RAND_1585[31:0];
  _RAND_1586 = {1{`RANDOM}};
  reg_csr_1586 = _RAND_1586[31:0];
  _RAND_1587 = {1{`RANDOM}};
  reg_csr_1587 = _RAND_1587[31:0];
  _RAND_1588 = {1{`RANDOM}};
  reg_csr_1588 = _RAND_1588[31:0];
  _RAND_1589 = {1{`RANDOM}};
  reg_csr_1589 = _RAND_1589[31:0];
  _RAND_1590 = {1{`RANDOM}};
  reg_csr_1590 = _RAND_1590[31:0];
  _RAND_1591 = {1{`RANDOM}};
  reg_csr_1591 = _RAND_1591[31:0];
  _RAND_1592 = {1{`RANDOM}};
  reg_csr_1592 = _RAND_1592[31:0];
  _RAND_1593 = {1{`RANDOM}};
  reg_csr_1593 = _RAND_1593[31:0];
  _RAND_1594 = {1{`RANDOM}};
  reg_csr_1594 = _RAND_1594[31:0];
  _RAND_1595 = {1{`RANDOM}};
  reg_csr_1595 = _RAND_1595[31:0];
  _RAND_1596 = {1{`RANDOM}};
  reg_csr_1596 = _RAND_1596[31:0];
  _RAND_1597 = {1{`RANDOM}};
  reg_csr_1597 = _RAND_1597[31:0];
  _RAND_1598 = {1{`RANDOM}};
  reg_csr_1598 = _RAND_1598[31:0];
  _RAND_1599 = {1{`RANDOM}};
  reg_csr_1599 = _RAND_1599[31:0];
  _RAND_1600 = {1{`RANDOM}};
  reg_csr_1600 = _RAND_1600[31:0];
  _RAND_1601 = {1{`RANDOM}};
  reg_csr_1601 = _RAND_1601[31:0];
  _RAND_1602 = {1{`RANDOM}};
  reg_csr_1602 = _RAND_1602[31:0];
  _RAND_1603 = {1{`RANDOM}};
  reg_csr_1603 = _RAND_1603[31:0];
  _RAND_1604 = {1{`RANDOM}};
  reg_csr_1604 = _RAND_1604[31:0];
  _RAND_1605 = {1{`RANDOM}};
  reg_csr_1605 = _RAND_1605[31:0];
  _RAND_1606 = {1{`RANDOM}};
  reg_csr_1606 = _RAND_1606[31:0];
  _RAND_1607 = {1{`RANDOM}};
  reg_csr_1607 = _RAND_1607[31:0];
  _RAND_1608 = {1{`RANDOM}};
  reg_csr_1608 = _RAND_1608[31:0];
  _RAND_1609 = {1{`RANDOM}};
  reg_csr_1609 = _RAND_1609[31:0];
  _RAND_1610 = {1{`RANDOM}};
  reg_csr_1610 = _RAND_1610[31:0];
  _RAND_1611 = {1{`RANDOM}};
  reg_csr_1611 = _RAND_1611[31:0];
  _RAND_1612 = {1{`RANDOM}};
  reg_csr_1612 = _RAND_1612[31:0];
  _RAND_1613 = {1{`RANDOM}};
  reg_csr_1613 = _RAND_1613[31:0];
  _RAND_1614 = {1{`RANDOM}};
  reg_csr_1614 = _RAND_1614[31:0];
  _RAND_1615 = {1{`RANDOM}};
  reg_csr_1615 = _RAND_1615[31:0];
  _RAND_1616 = {1{`RANDOM}};
  reg_csr_1616 = _RAND_1616[31:0];
  _RAND_1617 = {1{`RANDOM}};
  reg_csr_1617 = _RAND_1617[31:0];
  _RAND_1618 = {1{`RANDOM}};
  reg_csr_1618 = _RAND_1618[31:0];
  _RAND_1619 = {1{`RANDOM}};
  reg_csr_1619 = _RAND_1619[31:0];
  _RAND_1620 = {1{`RANDOM}};
  reg_csr_1620 = _RAND_1620[31:0];
  _RAND_1621 = {1{`RANDOM}};
  reg_csr_1621 = _RAND_1621[31:0];
  _RAND_1622 = {1{`RANDOM}};
  reg_csr_1622 = _RAND_1622[31:0];
  _RAND_1623 = {1{`RANDOM}};
  reg_csr_1623 = _RAND_1623[31:0];
  _RAND_1624 = {1{`RANDOM}};
  reg_csr_1624 = _RAND_1624[31:0];
  _RAND_1625 = {1{`RANDOM}};
  reg_csr_1625 = _RAND_1625[31:0];
  _RAND_1626 = {1{`RANDOM}};
  reg_csr_1626 = _RAND_1626[31:0];
  _RAND_1627 = {1{`RANDOM}};
  reg_csr_1627 = _RAND_1627[31:0];
  _RAND_1628 = {1{`RANDOM}};
  reg_csr_1628 = _RAND_1628[31:0];
  _RAND_1629 = {1{`RANDOM}};
  reg_csr_1629 = _RAND_1629[31:0];
  _RAND_1630 = {1{`RANDOM}};
  reg_csr_1630 = _RAND_1630[31:0];
  _RAND_1631 = {1{`RANDOM}};
  reg_csr_1631 = _RAND_1631[31:0];
  _RAND_1632 = {1{`RANDOM}};
  reg_csr_1632 = _RAND_1632[31:0];
  _RAND_1633 = {1{`RANDOM}};
  reg_csr_1633 = _RAND_1633[31:0];
  _RAND_1634 = {1{`RANDOM}};
  reg_csr_1634 = _RAND_1634[31:0];
  _RAND_1635 = {1{`RANDOM}};
  reg_csr_1635 = _RAND_1635[31:0];
  _RAND_1636 = {1{`RANDOM}};
  reg_csr_1636 = _RAND_1636[31:0];
  _RAND_1637 = {1{`RANDOM}};
  reg_csr_1637 = _RAND_1637[31:0];
  _RAND_1638 = {1{`RANDOM}};
  reg_csr_1638 = _RAND_1638[31:0];
  _RAND_1639 = {1{`RANDOM}};
  reg_csr_1639 = _RAND_1639[31:0];
  _RAND_1640 = {1{`RANDOM}};
  reg_csr_1640 = _RAND_1640[31:0];
  _RAND_1641 = {1{`RANDOM}};
  reg_csr_1641 = _RAND_1641[31:0];
  _RAND_1642 = {1{`RANDOM}};
  reg_csr_1642 = _RAND_1642[31:0];
  _RAND_1643 = {1{`RANDOM}};
  reg_csr_1643 = _RAND_1643[31:0];
  _RAND_1644 = {1{`RANDOM}};
  reg_csr_1644 = _RAND_1644[31:0];
  _RAND_1645 = {1{`RANDOM}};
  reg_csr_1645 = _RAND_1645[31:0];
  _RAND_1646 = {1{`RANDOM}};
  reg_csr_1646 = _RAND_1646[31:0];
  _RAND_1647 = {1{`RANDOM}};
  reg_csr_1647 = _RAND_1647[31:0];
  _RAND_1648 = {1{`RANDOM}};
  reg_csr_1648 = _RAND_1648[31:0];
  _RAND_1649 = {1{`RANDOM}};
  reg_csr_1649 = _RAND_1649[31:0];
  _RAND_1650 = {1{`RANDOM}};
  reg_csr_1650 = _RAND_1650[31:0];
  _RAND_1651 = {1{`RANDOM}};
  reg_csr_1651 = _RAND_1651[31:0];
  _RAND_1652 = {1{`RANDOM}};
  reg_csr_1652 = _RAND_1652[31:0];
  _RAND_1653 = {1{`RANDOM}};
  reg_csr_1653 = _RAND_1653[31:0];
  _RAND_1654 = {1{`RANDOM}};
  reg_csr_1654 = _RAND_1654[31:0];
  _RAND_1655 = {1{`RANDOM}};
  reg_csr_1655 = _RAND_1655[31:0];
  _RAND_1656 = {1{`RANDOM}};
  reg_csr_1656 = _RAND_1656[31:0];
  _RAND_1657 = {1{`RANDOM}};
  reg_csr_1657 = _RAND_1657[31:0];
  _RAND_1658 = {1{`RANDOM}};
  reg_csr_1658 = _RAND_1658[31:0];
  _RAND_1659 = {1{`RANDOM}};
  reg_csr_1659 = _RAND_1659[31:0];
  _RAND_1660 = {1{`RANDOM}};
  reg_csr_1660 = _RAND_1660[31:0];
  _RAND_1661 = {1{`RANDOM}};
  reg_csr_1661 = _RAND_1661[31:0];
  _RAND_1662 = {1{`RANDOM}};
  reg_csr_1662 = _RAND_1662[31:0];
  _RAND_1663 = {1{`RANDOM}};
  reg_csr_1663 = _RAND_1663[31:0];
  _RAND_1664 = {1{`RANDOM}};
  reg_csr_1664 = _RAND_1664[31:0];
  _RAND_1665 = {1{`RANDOM}};
  reg_csr_1665 = _RAND_1665[31:0];
  _RAND_1666 = {1{`RANDOM}};
  reg_csr_1666 = _RAND_1666[31:0];
  _RAND_1667 = {1{`RANDOM}};
  reg_csr_1667 = _RAND_1667[31:0];
  _RAND_1668 = {1{`RANDOM}};
  reg_csr_1668 = _RAND_1668[31:0];
  _RAND_1669 = {1{`RANDOM}};
  reg_csr_1669 = _RAND_1669[31:0];
  _RAND_1670 = {1{`RANDOM}};
  reg_csr_1670 = _RAND_1670[31:0];
  _RAND_1671 = {1{`RANDOM}};
  reg_csr_1671 = _RAND_1671[31:0];
  _RAND_1672 = {1{`RANDOM}};
  reg_csr_1672 = _RAND_1672[31:0];
  _RAND_1673 = {1{`RANDOM}};
  reg_csr_1673 = _RAND_1673[31:0];
  _RAND_1674 = {1{`RANDOM}};
  reg_csr_1674 = _RAND_1674[31:0];
  _RAND_1675 = {1{`RANDOM}};
  reg_csr_1675 = _RAND_1675[31:0];
  _RAND_1676 = {1{`RANDOM}};
  reg_csr_1676 = _RAND_1676[31:0];
  _RAND_1677 = {1{`RANDOM}};
  reg_csr_1677 = _RAND_1677[31:0];
  _RAND_1678 = {1{`RANDOM}};
  reg_csr_1678 = _RAND_1678[31:0];
  _RAND_1679 = {1{`RANDOM}};
  reg_csr_1679 = _RAND_1679[31:0];
  _RAND_1680 = {1{`RANDOM}};
  reg_csr_1680 = _RAND_1680[31:0];
  _RAND_1681 = {1{`RANDOM}};
  reg_csr_1681 = _RAND_1681[31:0];
  _RAND_1682 = {1{`RANDOM}};
  reg_csr_1682 = _RAND_1682[31:0];
  _RAND_1683 = {1{`RANDOM}};
  reg_csr_1683 = _RAND_1683[31:0];
  _RAND_1684 = {1{`RANDOM}};
  reg_csr_1684 = _RAND_1684[31:0];
  _RAND_1685 = {1{`RANDOM}};
  reg_csr_1685 = _RAND_1685[31:0];
  _RAND_1686 = {1{`RANDOM}};
  reg_csr_1686 = _RAND_1686[31:0];
  _RAND_1687 = {1{`RANDOM}};
  reg_csr_1687 = _RAND_1687[31:0];
  _RAND_1688 = {1{`RANDOM}};
  reg_csr_1688 = _RAND_1688[31:0];
  _RAND_1689 = {1{`RANDOM}};
  reg_csr_1689 = _RAND_1689[31:0];
  _RAND_1690 = {1{`RANDOM}};
  reg_csr_1690 = _RAND_1690[31:0];
  _RAND_1691 = {1{`RANDOM}};
  reg_csr_1691 = _RAND_1691[31:0];
  _RAND_1692 = {1{`RANDOM}};
  reg_csr_1692 = _RAND_1692[31:0];
  _RAND_1693 = {1{`RANDOM}};
  reg_csr_1693 = _RAND_1693[31:0];
  _RAND_1694 = {1{`RANDOM}};
  reg_csr_1694 = _RAND_1694[31:0];
  _RAND_1695 = {1{`RANDOM}};
  reg_csr_1695 = _RAND_1695[31:0];
  _RAND_1696 = {1{`RANDOM}};
  reg_csr_1696 = _RAND_1696[31:0];
  _RAND_1697 = {1{`RANDOM}};
  reg_csr_1697 = _RAND_1697[31:0];
  _RAND_1698 = {1{`RANDOM}};
  reg_csr_1698 = _RAND_1698[31:0];
  _RAND_1699 = {1{`RANDOM}};
  reg_csr_1699 = _RAND_1699[31:0];
  _RAND_1700 = {1{`RANDOM}};
  reg_csr_1700 = _RAND_1700[31:0];
  _RAND_1701 = {1{`RANDOM}};
  reg_csr_1701 = _RAND_1701[31:0];
  _RAND_1702 = {1{`RANDOM}};
  reg_csr_1702 = _RAND_1702[31:0];
  _RAND_1703 = {1{`RANDOM}};
  reg_csr_1703 = _RAND_1703[31:0];
  _RAND_1704 = {1{`RANDOM}};
  reg_csr_1704 = _RAND_1704[31:0];
  _RAND_1705 = {1{`RANDOM}};
  reg_csr_1705 = _RAND_1705[31:0];
  _RAND_1706 = {1{`RANDOM}};
  reg_csr_1706 = _RAND_1706[31:0];
  _RAND_1707 = {1{`RANDOM}};
  reg_csr_1707 = _RAND_1707[31:0];
  _RAND_1708 = {1{`RANDOM}};
  reg_csr_1708 = _RAND_1708[31:0];
  _RAND_1709 = {1{`RANDOM}};
  reg_csr_1709 = _RAND_1709[31:0];
  _RAND_1710 = {1{`RANDOM}};
  reg_csr_1710 = _RAND_1710[31:0];
  _RAND_1711 = {1{`RANDOM}};
  reg_csr_1711 = _RAND_1711[31:0];
  _RAND_1712 = {1{`RANDOM}};
  reg_csr_1712 = _RAND_1712[31:0];
  _RAND_1713 = {1{`RANDOM}};
  reg_csr_1713 = _RAND_1713[31:0];
  _RAND_1714 = {1{`RANDOM}};
  reg_csr_1714 = _RAND_1714[31:0];
  _RAND_1715 = {1{`RANDOM}};
  reg_csr_1715 = _RAND_1715[31:0];
  _RAND_1716 = {1{`RANDOM}};
  reg_csr_1716 = _RAND_1716[31:0];
  _RAND_1717 = {1{`RANDOM}};
  reg_csr_1717 = _RAND_1717[31:0];
  _RAND_1718 = {1{`RANDOM}};
  reg_csr_1718 = _RAND_1718[31:0];
  _RAND_1719 = {1{`RANDOM}};
  reg_csr_1719 = _RAND_1719[31:0];
  _RAND_1720 = {1{`RANDOM}};
  reg_csr_1720 = _RAND_1720[31:0];
  _RAND_1721 = {1{`RANDOM}};
  reg_csr_1721 = _RAND_1721[31:0];
  _RAND_1722 = {1{`RANDOM}};
  reg_csr_1722 = _RAND_1722[31:0];
  _RAND_1723 = {1{`RANDOM}};
  reg_csr_1723 = _RAND_1723[31:0];
  _RAND_1724 = {1{`RANDOM}};
  reg_csr_1724 = _RAND_1724[31:0];
  _RAND_1725 = {1{`RANDOM}};
  reg_csr_1725 = _RAND_1725[31:0];
  _RAND_1726 = {1{`RANDOM}};
  reg_csr_1726 = _RAND_1726[31:0];
  _RAND_1727 = {1{`RANDOM}};
  reg_csr_1727 = _RAND_1727[31:0];
  _RAND_1728 = {1{`RANDOM}};
  reg_csr_1728 = _RAND_1728[31:0];
  _RAND_1729 = {1{`RANDOM}};
  reg_csr_1729 = _RAND_1729[31:0];
  _RAND_1730 = {1{`RANDOM}};
  reg_csr_1730 = _RAND_1730[31:0];
  _RAND_1731 = {1{`RANDOM}};
  reg_csr_1731 = _RAND_1731[31:0];
  _RAND_1732 = {1{`RANDOM}};
  reg_csr_1732 = _RAND_1732[31:0];
  _RAND_1733 = {1{`RANDOM}};
  reg_csr_1733 = _RAND_1733[31:0];
  _RAND_1734 = {1{`RANDOM}};
  reg_csr_1734 = _RAND_1734[31:0];
  _RAND_1735 = {1{`RANDOM}};
  reg_csr_1735 = _RAND_1735[31:0];
  _RAND_1736 = {1{`RANDOM}};
  reg_csr_1736 = _RAND_1736[31:0];
  _RAND_1737 = {1{`RANDOM}};
  reg_csr_1737 = _RAND_1737[31:0];
  _RAND_1738 = {1{`RANDOM}};
  reg_csr_1738 = _RAND_1738[31:0];
  _RAND_1739 = {1{`RANDOM}};
  reg_csr_1739 = _RAND_1739[31:0];
  _RAND_1740 = {1{`RANDOM}};
  reg_csr_1740 = _RAND_1740[31:0];
  _RAND_1741 = {1{`RANDOM}};
  reg_csr_1741 = _RAND_1741[31:0];
  _RAND_1742 = {1{`RANDOM}};
  reg_csr_1742 = _RAND_1742[31:0];
  _RAND_1743 = {1{`RANDOM}};
  reg_csr_1743 = _RAND_1743[31:0];
  _RAND_1744 = {1{`RANDOM}};
  reg_csr_1744 = _RAND_1744[31:0];
  _RAND_1745 = {1{`RANDOM}};
  reg_csr_1745 = _RAND_1745[31:0];
  _RAND_1746 = {1{`RANDOM}};
  reg_csr_1746 = _RAND_1746[31:0];
  _RAND_1747 = {1{`RANDOM}};
  reg_csr_1747 = _RAND_1747[31:0];
  _RAND_1748 = {1{`RANDOM}};
  reg_csr_1748 = _RAND_1748[31:0];
  _RAND_1749 = {1{`RANDOM}};
  reg_csr_1749 = _RAND_1749[31:0];
  _RAND_1750 = {1{`RANDOM}};
  reg_csr_1750 = _RAND_1750[31:0];
  _RAND_1751 = {1{`RANDOM}};
  reg_csr_1751 = _RAND_1751[31:0];
  _RAND_1752 = {1{`RANDOM}};
  reg_csr_1752 = _RAND_1752[31:0];
  _RAND_1753 = {1{`RANDOM}};
  reg_csr_1753 = _RAND_1753[31:0];
  _RAND_1754 = {1{`RANDOM}};
  reg_csr_1754 = _RAND_1754[31:0];
  _RAND_1755 = {1{`RANDOM}};
  reg_csr_1755 = _RAND_1755[31:0];
  _RAND_1756 = {1{`RANDOM}};
  reg_csr_1756 = _RAND_1756[31:0];
  _RAND_1757 = {1{`RANDOM}};
  reg_csr_1757 = _RAND_1757[31:0];
  _RAND_1758 = {1{`RANDOM}};
  reg_csr_1758 = _RAND_1758[31:0];
  _RAND_1759 = {1{`RANDOM}};
  reg_csr_1759 = _RAND_1759[31:0];
  _RAND_1760 = {1{`RANDOM}};
  reg_csr_1760 = _RAND_1760[31:0];
  _RAND_1761 = {1{`RANDOM}};
  reg_csr_1761 = _RAND_1761[31:0];
  _RAND_1762 = {1{`RANDOM}};
  reg_csr_1762 = _RAND_1762[31:0];
  _RAND_1763 = {1{`RANDOM}};
  reg_csr_1763 = _RAND_1763[31:0];
  _RAND_1764 = {1{`RANDOM}};
  reg_csr_1764 = _RAND_1764[31:0];
  _RAND_1765 = {1{`RANDOM}};
  reg_csr_1765 = _RAND_1765[31:0];
  _RAND_1766 = {1{`RANDOM}};
  reg_csr_1766 = _RAND_1766[31:0];
  _RAND_1767 = {1{`RANDOM}};
  reg_csr_1767 = _RAND_1767[31:0];
  _RAND_1768 = {1{`RANDOM}};
  reg_csr_1768 = _RAND_1768[31:0];
  _RAND_1769 = {1{`RANDOM}};
  reg_csr_1769 = _RAND_1769[31:0];
  _RAND_1770 = {1{`RANDOM}};
  reg_csr_1770 = _RAND_1770[31:0];
  _RAND_1771 = {1{`RANDOM}};
  reg_csr_1771 = _RAND_1771[31:0];
  _RAND_1772 = {1{`RANDOM}};
  reg_csr_1772 = _RAND_1772[31:0];
  _RAND_1773 = {1{`RANDOM}};
  reg_csr_1773 = _RAND_1773[31:0];
  _RAND_1774 = {1{`RANDOM}};
  reg_csr_1774 = _RAND_1774[31:0];
  _RAND_1775 = {1{`RANDOM}};
  reg_csr_1775 = _RAND_1775[31:0];
  _RAND_1776 = {1{`RANDOM}};
  reg_csr_1776 = _RAND_1776[31:0];
  _RAND_1777 = {1{`RANDOM}};
  reg_csr_1777 = _RAND_1777[31:0];
  _RAND_1778 = {1{`RANDOM}};
  reg_csr_1778 = _RAND_1778[31:0];
  _RAND_1779 = {1{`RANDOM}};
  reg_csr_1779 = _RAND_1779[31:0];
  _RAND_1780 = {1{`RANDOM}};
  reg_csr_1780 = _RAND_1780[31:0];
  _RAND_1781 = {1{`RANDOM}};
  reg_csr_1781 = _RAND_1781[31:0];
  _RAND_1782 = {1{`RANDOM}};
  reg_csr_1782 = _RAND_1782[31:0];
  _RAND_1783 = {1{`RANDOM}};
  reg_csr_1783 = _RAND_1783[31:0];
  _RAND_1784 = {1{`RANDOM}};
  reg_csr_1784 = _RAND_1784[31:0];
  _RAND_1785 = {1{`RANDOM}};
  reg_csr_1785 = _RAND_1785[31:0];
  _RAND_1786 = {1{`RANDOM}};
  reg_csr_1786 = _RAND_1786[31:0];
  _RAND_1787 = {1{`RANDOM}};
  reg_csr_1787 = _RAND_1787[31:0];
  _RAND_1788 = {1{`RANDOM}};
  reg_csr_1788 = _RAND_1788[31:0];
  _RAND_1789 = {1{`RANDOM}};
  reg_csr_1789 = _RAND_1789[31:0];
  _RAND_1790 = {1{`RANDOM}};
  reg_csr_1790 = _RAND_1790[31:0];
  _RAND_1791 = {1{`RANDOM}};
  reg_csr_1791 = _RAND_1791[31:0];
  _RAND_1792 = {1{`RANDOM}};
  reg_csr_1792 = _RAND_1792[31:0];
  _RAND_1793 = {1{`RANDOM}};
  reg_csr_1793 = _RAND_1793[31:0];
  _RAND_1794 = {1{`RANDOM}};
  reg_csr_1794 = _RAND_1794[31:0];
  _RAND_1795 = {1{`RANDOM}};
  reg_csr_1795 = _RAND_1795[31:0];
  _RAND_1796 = {1{`RANDOM}};
  reg_csr_1796 = _RAND_1796[31:0];
  _RAND_1797 = {1{`RANDOM}};
  reg_csr_1797 = _RAND_1797[31:0];
  _RAND_1798 = {1{`RANDOM}};
  reg_csr_1798 = _RAND_1798[31:0];
  _RAND_1799 = {1{`RANDOM}};
  reg_csr_1799 = _RAND_1799[31:0];
  _RAND_1800 = {1{`RANDOM}};
  reg_csr_1800 = _RAND_1800[31:0];
  _RAND_1801 = {1{`RANDOM}};
  reg_csr_1801 = _RAND_1801[31:0];
  _RAND_1802 = {1{`RANDOM}};
  reg_csr_1802 = _RAND_1802[31:0];
  _RAND_1803 = {1{`RANDOM}};
  reg_csr_1803 = _RAND_1803[31:0];
  _RAND_1804 = {1{`RANDOM}};
  reg_csr_1804 = _RAND_1804[31:0];
  _RAND_1805 = {1{`RANDOM}};
  reg_csr_1805 = _RAND_1805[31:0];
  _RAND_1806 = {1{`RANDOM}};
  reg_csr_1806 = _RAND_1806[31:0];
  _RAND_1807 = {1{`RANDOM}};
  reg_csr_1807 = _RAND_1807[31:0];
  _RAND_1808 = {1{`RANDOM}};
  reg_csr_1808 = _RAND_1808[31:0];
  _RAND_1809 = {1{`RANDOM}};
  reg_csr_1809 = _RAND_1809[31:0];
  _RAND_1810 = {1{`RANDOM}};
  reg_csr_1810 = _RAND_1810[31:0];
  _RAND_1811 = {1{`RANDOM}};
  reg_csr_1811 = _RAND_1811[31:0];
  _RAND_1812 = {1{`RANDOM}};
  reg_csr_1812 = _RAND_1812[31:0];
  _RAND_1813 = {1{`RANDOM}};
  reg_csr_1813 = _RAND_1813[31:0];
  _RAND_1814 = {1{`RANDOM}};
  reg_csr_1814 = _RAND_1814[31:0];
  _RAND_1815 = {1{`RANDOM}};
  reg_csr_1815 = _RAND_1815[31:0];
  _RAND_1816 = {1{`RANDOM}};
  reg_csr_1816 = _RAND_1816[31:0];
  _RAND_1817 = {1{`RANDOM}};
  reg_csr_1817 = _RAND_1817[31:0];
  _RAND_1818 = {1{`RANDOM}};
  reg_csr_1818 = _RAND_1818[31:0];
  _RAND_1819 = {1{`RANDOM}};
  reg_csr_1819 = _RAND_1819[31:0];
  _RAND_1820 = {1{`RANDOM}};
  reg_csr_1820 = _RAND_1820[31:0];
  _RAND_1821 = {1{`RANDOM}};
  reg_csr_1821 = _RAND_1821[31:0];
  _RAND_1822 = {1{`RANDOM}};
  reg_csr_1822 = _RAND_1822[31:0];
  _RAND_1823 = {1{`RANDOM}};
  reg_csr_1823 = _RAND_1823[31:0];
  _RAND_1824 = {1{`RANDOM}};
  reg_csr_1824 = _RAND_1824[31:0];
  _RAND_1825 = {1{`RANDOM}};
  reg_csr_1825 = _RAND_1825[31:0];
  _RAND_1826 = {1{`RANDOM}};
  reg_csr_1826 = _RAND_1826[31:0];
  _RAND_1827 = {1{`RANDOM}};
  reg_csr_1827 = _RAND_1827[31:0];
  _RAND_1828 = {1{`RANDOM}};
  reg_csr_1828 = _RAND_1828[31:0];
  _RAND_1829 = {1{`RANDOM}};
  reg_csr_1829 = _RAND_1829[31:0];
  _RAND_1830 = {1{`RANDOM}};
  reg_csr_1830 = _RAND_1830[31:0];
  _RAND_1831 = {1{`RANDOM}};
  reg_csr_1831 = _RAND_1831[31:0];
  _RAND_1832 = {1{`RANDOM}};
  reg_csr_1832 = _RAND_1832[31:0];
  _RAND_1833 = {1{`RANDOM}};
  reg_csr_1833 = _RAND_1833[31:0];
  _RAND_1834 = {1{`RANDOM}};
  reg_csr_1834 = _RAND_1834[31:0];
  _RAND_1835 = {1{`RANDOM}};
  reg_csr_1835 = _RAND_1835[31:0];
  _RAND_1836 = {1{`RANDOM}};
  reg_csr_1836 = _RAND_1836[31:0];
  _RAND_1837 = {1{`RANDOM}};
  reg_csr_1837 = _RAND_1837[31:0];
  _RAND_1838 = {1{`RANDOM}};
  reg_csr_1838 = _RAND_1838[31:0];
  _RAND_1839 = {1{`RANDOM}};
  reg_csr_1839 = _RAND_1839[31:0];
  _RAND_1840 = {1{`RANDOM}};
  reg_csr_1840 = _RAND_1840[31:0];
  _RAND_1841 = {1{`RANDOM}};
  reg_csr_1841 = _RAND_1841[31:0];
  _RAND_1842 = {1{`RANDOM}};
  reg_csr_1842 = _RAND_1842[31:0];
  _RAND_1843 = {1{`RANDOM}};
  reg_csr_1843 = _RAND_1843[31:0];
  _RAND_1844 = {1{`RANDOM}};
  reg_csr_1844 = _RAND_1844[31:0];
  _RAND_1845 = {1{`RANDOM}};
  reg_csr_1845 = _RAND_1845[31:0];
  _RAND_1846 = {1{`RANDOM}};
  reg_csr_1846 = _RAND_1846[31:0];
  _RAND_1847 = {1{`RANDOM}};
  reg_csr_1847 = _RAND_1847[31:0];
  _RAND_1848 = {1{`RANDOM}};
  reg_csr_1848 = _RAND_1848[31:0];
  _RAND_1849 = {1{`RANDOM}};
  reg_csr_1849 = _RAND_1849[31:0];
  _RAND_1850 = {1{`RANDOM}};
  reg_csr_1850 = _RAND_1850[31:0];
  _RAND_1851 = {1{`RANDOM}};
  reg_csr_1851 = _RAND_1851[31:0];
  _RAND_1852 = {1{`RANDOM}};
  reg_csr_1852 = _RAND_1852[31:0];
  _RAND_1853 = {1{`RANDOM}};
  reg_csr_1853 = _RAND_1853[31:0];
  _RAND_1854 = {1{`RANDOM}};
  reg_csr_1854 = _RAND_1854[31:0];
  _RAND_1855 = {1{`RANDOM}};
  reg_csr_1855 = _RAND_1855[31:0];
  _RAND_1856 = {1{`RANDOM}};
  reg_csr_1856 = _RAND_1856[31:0];
  _RAND_1857 = {1{`RANDOM}};
  reg_csr_1857 = _RAND_1857[31:0];
  _RAND_1858 = {1{`RANDOM}};
  reg_csr_1858 = _RAND_1858[31:0];
  _RAND_1859 = {1{`RANDOM}};
  reg_csr_1859 = _RAND_1859[31:0];
  _RAND_1860 = {1{`RANDOM}};
  reg_csr_1860 = _RAND_1860[31:0];
  _RAND_1861 = {1{`RANDOM}};
  reg_csr_1861 = _RAND_1861[31:0];
  _RAND_1862 = {1{`RANDOM}};
  reg_csr_1862 = _RAND_1862[31:0];
  _RAND_1863 = {1{`RANDOM}};
  reg_csr_1863 = _RAND_1863[31:0];
  _RAND_1864 = {1{`RANDOM}};
  reg_csr_1864 = _RAND_1864[31:0];
  _RAND_1865 = {1{`RANDOM}};
  reg_csr_1865 = _RAND_1865[31:0];
  _RAND_1866 = {1{`RANDOM}};
  reg_csr_1866 = _RAND_1866[31:0];
  _RAND_1867 = {1{`RANDOM}};
  reg_csr_1867 = _RAND_1867[31:0];
  _RAND_1868 = {1{`RANDOM}};
  reg_csr_1868 = _RAND_1868[31:0];
  _RAND_1869 = {1{`RANDOM}};
  reg_csr_1869 = _RAND_1869[31:0];
  _RAND_1870 = {1{`RANDOM}};
  reg_csr_1870 = _RAND_1870[31:0];
  _RAND_1871 = {1{`RANDOM}};
  reg_csr_1871 = _RAND_1871[31:0];
  _RAND_1872 = {1{`RANDOM}};
  reg_csr_1872 = _RAND_1872[31:0];
  _RAND_1873 = {1{`RANDOM}};
  reg_csr_1873 = _RAND_1873[31:0];
  _RAND_1874 = {1{`RANDOM}};
  reg_csr_1874 = _RAND_1874[31:0];
  _RAND_1875 = {1{`RANDOM}};
  reg_csr_1875 = _RAND_1875[31:0];
  _RAND_1876 = {1{`RANDOM}};
  reg_csr_1876 = _RAND_1876[31:0];
  _RAND_1877 = {1{`RANDOM}};
  reg_csr_1877 = _RAND_1877[31:0];
  _RAND_1878 = {1{`RANDOM}};
  reg_csr_1878 = _RAND_1878[31:0];
  _RAND_1879 = {1{`RANDOM}};
  reg_csr_1879 = _RAND_1879[31:0];
  _RAND_1880 = {1{`RANDOM}};
  reg_csr_1880 = _RAND_1880[31:0];
  _RAND_1881 = {1{`RANDOM}};
  reg_csr_1881 = _RAND_1881[31:0];
  _RAND_1882 = {1{`RANDOM}};
  reg_csr_1882 = _RAND_1882[31:0];
  _RAND_1883 = {1{`RANDOM}};
  reg_csr_1883 = _RAND_1883[31:0];
  _RAND_1884 = {1{`RANDOM}};
  reg_csr_1884 = _RAND_1884[31:0];
  _RAND_1885 = {1{`RANDOM}};
  reg_csr_1885 = _RAND_1885[31:0];
  _RAND_1886 = {1{`RANDOM}};
  reg_csr_1886 = _RAND_1886[31:0];
  _RAND_1887 = {1{`RANDOM}};
  reg_csr_1887 = _RAND_1887[31:0];
  _RAND_1888 = {1{`RANDOM}};
  reg_csr_1888 = _RAND_1888[31:0];
  _RAND_1889 = {1{`RANDOM}};
  reg_csr_1889 = _RAND_1889[31:0];
  _RAND_1890 = {1{`RANDOM}};
  reg_csr_1890 = _RAND_1890[31:0];
  _RAND_1891 = {1{`RANDOM}};
  reg_csr_1891 = _RAND_1891[31:0];
  _RAND_1892 = {1{`RANDOM}};
  reg_csr_1892 = _RAND_1892[31:0];
  _RAND_1893 = {1{`RANDOM}};
  reg_csr_1893 = _RAND_1893[31:0];
  _RAND_1894 = {1{`RANDOM}};
  reg_csr_1894 = _RAND_1894[31:0];
  _RAND_1895 = {1{`RANDOM}};
  reg_csr_1895 = _RAND_1895[31:0];
  _RAND_1896 = {1{`RANDOM}};
  reg_csr_1896 = _RAND_1896[31:0];
  _RAND_1897 = {1{`RANDOM}};
  reg_csr_1897 = _RAND_1897[31:0];
  _RAND_1898 = {1{`RANDOM}};
  reg_csr_1898 = _RAND_1898[31:0];
  _RAND_1899 = {1{`RANDOM}};
  reg_csr_1899 = _RAND_1899[31:0];
  _RAND_1900 = {1{`RANDOM}};
  reg_csr_1900 = _RAND_1900[31:0];
  _RAND_1901 = {1{`RANDOM}};
  reg_csr_1901 = _RAND_1901[31:0];
  _RAND_1902 = {1{`RANDOM}};
  reg_csr_1902 = _RAND_1902[31:0];
  _RAND_1903 = {1{`RANDOM}};
  reg_csr_1903 = _RAND_1903[31:0];
  _RAND_1904 = {1{`RANDOM}};
  reg_csr_1904 = _RAND_1904[31:0];
  _RAND_1905 = {1{`RANDOM}};
  reg_csr_1905 = _RAND_1905[31:0];
  _RAND_1906 = {1{`RANDOM}};
  reg_csr_1906 = _RAND_1906[31:0];
  _RAND_1907 = {1{`RANDOM}};
  reg_csr_1907 = _RAND_1907[31:0];
  _RAND_1908 = {1{`RANDOM}};
  reg_csr_1908 = _RAND_1908[31:0];
  _RAND_1909 = {1{`RANDOM}};
  reg_csr_1909 = _RAND_1909[31:0];
  _RAND_1910 = {1{`RANDOM}};
  reg_csr_1910 = _RAND_1910[31:0];
  _RAND_1911 = {1{`RANDOM}};
  reg_csr_1911 = _RAND_1911[31:0];
  _RAND_1912 = {1{`RANDOM}};
  reg_csr_1912 = _RAND_1912[31:0];
  _RAND_1913 = {1{`RANDOM}};
  reg_csr_1913 = _RAND_1913[31:0];
  _RAND_1914 = {1{`RANDOM}};
  reg_csr_1914 = _RAND_1914[31:0];
  _RAND_1915 = {1{`RANDOM}};
  reg_csr_1915 = _RAND_1915[31:0];
  _RAND_1916 = {1{`RANDOM}};
  reg_csr_1916 = _RAND_1916[31:0];
  _RAND_1917 = {1{`RANDOM}};
  reg_csr_1917 = _RAND_1917[31:0];
  _RAND_1918 = {1{`RANDOM}};
  reg_csr_1918 = _RAND_1918[31:0];
  _RAND_1919 = {1{`RANDOM}};
  reg_csr_1919 = _RAND_1919[31:0];
  _RAND_1920 = {1{`RANDOM}};
  reg_csr_1920 = _RAND_1920[31:0];
  _RAND_1921 = {1{`RANDOM}};
  reg_csr_1921 = _RAND_1921[31:0];
  _RAND_1922 = {1{`RANDOM}};
  reg_csr_1922 = _RAND_1922[31:0];
  _RAND_1923 = {1{`RANDOM}};
  reg_csr_1923 = _RAND_1923[31:0];
  _RAND_1924 = {1{`RANDOM}};
  reg_csr_1924 = _RAND_1924[31:0];
  _RAND_1925 = {1{`RANDOM}};
  reg_csr_1925 = _RAND_1925[31:0];
  _RAND_1926 = {1{`RANDOM}};
  reg_csr_1926 = _RAND_1926[31:0];
  _RAND_1927 = {1{`RANDOM}};
  reg_csr_1927 = _RAND_1927[31:0];
  _RAND_1928 = {1{`RANDOM}};
  reg_csr_1928 = _RAND_1928[31:0];
  _RAND_1929 = {1{`RANDOM}};
  reg_csr_1929 = _RAND_1929[31:0];
  _RAND_1930 = {1{`RANDOM}};
  reg_csr_1930 = _RAND_1930[31:0];
  _RAND_1931 = {1{`RANDOM}};
  reg_csr_1931 = _RAND_1931[31:0];
  _RAND_1932 = {1{`RANDOM}};
  reg_csr_1932 = _RAND_1932[31:0];
  _RAND_1933 = {1{`RANDOM}};
  reg_csr_1933 = _RAND_1933[31:0];
  _RAND_1934 = {1{`RANDOM}};
  reg_csr_1934 = _RAND_1934[31:0];
  _RAND_1935 = {1{`RANDOM}};
  reg_csr_1935 = _RAND_1935[31:0];
  _RAND_1936 = {1{`RANDOM}};
  reg_csr_1936 = _RAND_1936[31:0];
  _RAND_1937 = {1{`RANDOM}};
  reg_csr_1937 = _RAND_1937[31:0];
  _RAND_1938 = {1{`RANDOM}};
  reg_csr_1938 = _RAND_1938[31:0];
  _RAND_1939 = {1{`RANDOM}};
  reg_csr_1939 = _RAND_1939[31:0];
  _RAND_1940 = {1{`RANDOM}};
  reg_csr_1940 = _RAND_1940[31:0];
  _RAND_1941 = {1{`RANDOM}};
  reg_csr_1941 = _RAND_1941[31:0];
  _RAND_1942 = {1{`RANDOM}};
  reg_csr_1942 = _RAND_1942[31:0];
  _RAND_1943 = {1{`RANDOM}};
  reg_csr_1943 = _RAND_1943[31:0];
  _RAND_1944 = {1{`RANDOM}};
  reg_csr_1944 = _RAND_1944[31:0];
  _RAND_1945 = {1{`RANDOM}};
  reg_csr_1945 = _RAND_1945[31:0];
  _RAND_1946 = {1{`RANDOM}};
  reg_csr_1946 = _RAND_1946[31:0];
  _RAND_1947 = {1{`RANDOM}};
  reg_csr_1947 = _RAND_1947[31:0];
  _RAND_1948 = {1{`RANDOM}};
  reg_csr_1948 = _RAND_1948[31:0];
  _RAND_1949 = {1{`RANDOM}};
  reg_csr_1949 = _RAND_1949[31:0];
  _RAND_1950 = {1{`RANDOM}};
  reg_csr_1950 = _RAND_1950[31:0];
  _RAND_1951 = {1{`RANDOM}};
  reg_csr_1951 = _RAND_1951[31:0];
  _RAND_1952 = {1{`RANDOM}};
  reg_csr_1952 = _RAND_1952[31:0];
  _RAND_1953 = {1{`RANDOM}};
  reg_csr_1953 = _RAND_1953[31:0];
  _RAND_1954 = {1{`RANDOM}};
  reg_csr_1954 = _RAND_1954[31:0];
  _RAND_1955 = {1{`RANDOM}};
  reg_csr_1955 = _RAND_1955[31:0];
  _RAND_1956 = {1{`RANDOM}};
  reg_csr_1956 = _RAND_1956[31:0];
  _RAND_1957 = {1{`RANDOM}};
  reg_csr_1957 = _RAND_1957[31:0];
  _RAND_1958 = {1{`RANDOM}};
  reg_csr_1958 = _RAND_1958[31:0];
  _RAND_1959 = {1{`RANDOM}};
  reg_csr_1959 = _RAND_1959[31:0];
  _RAND_1960 = {1{`RANDOM}};
  reg_csr_1960 = _RAND_1960[31:0];
  _RAND_1961 = {1{`RANDOM}};
  reg_csr_1961 = _RAND_1961[31:0];
  _RAND_1962 = {1{`RANDOM}};
  reg_csr_1962 = _RAND_1962[31:0];
  _RAND_1963 = {1{`RANDOM}};
  reg_csr_1963 = _RAND_1963[31:0];
  _RAND_1964 = {1{`RANDOM}};
  reg_csr_1964 = _RAND_1964[31:0];
  _RAND_1965 = {1{`RANDOM}};
  reg_csr_1965 = _RAND_1965[31:0];
  _RAND_1966 = {1{`RANDOM}};
  reg_csr_1966 = _RAND_1966[31:0];
  _RAND_1967 = {1{`RANDOM}};
  reg_csr_1967 = _RAND_1967[31:0];
  _RAND_1968 = {1{`RANDOM}};
  reg_csr_1968 = _RAND_1968[31:0];
  _RAND_1969 = {1{`RANDOM}};
  reg_csr_1969 = _RAND_1969[31:0];
  _RAND_1970 = {1{`RANDOM}};
  reg_csr_1970 = _RAND_1970[31:0];
  _RAND_1971 = {1{`RANDOM}};
  reg_csr_1971 = _RAND_1971[31:0];
  _RAND_1972 = {1{`RANDOM}};
  reg_csr_1972 = _RAND_1972[31:0];
  _RAND_1973 = {1{`RANDOM}};
  reg_csr_1973 = _RAND_1973[31:0];
  _RAND_1974 = {1{`RANDOM}};
  reg_csr_1974 = _RAND_1974[31:0];
  _RAND_1975 = {1{`RANDOM}};
  reg_csr_1975 = _RAND_1975[31:0];
  _RAND_1976 = {1{`RANDOM}};
  reg_csr_1976 = _RAND_1976[31:0];
  _RAND_1977 = {1{`RANDOM}};
  reg_csr_1977 = _RAND_1977[31:0];
  _RAND_1978 = {1{`RANDOM}};
  reg_csr_1978 = _RAND_1978[31:0];
  _RAND_1979 = {1{`RANDOM}};
  reg_csr_1979 = _RAND_1979[31:0];
  _RAND_1980 = {1{`RANDOM}};
  reg_csr_1980 = _RAND_1980[31:0];
  _RAND_1981 = {1{`RANDOM}};
  reg_csr_1981 = _RAND_1981[31:0];
  _RAND_1982 = {1{`RANDOM}};
  reg_csr_1982 = _RAND_1982[31:0];
  _RAND_1983 = {1{`RANDOM}};
  reg_csr_1983 = _RAND_1983[31:0];
  _RAND_1984 = {1{`RANDOM}};
  reg_csr_1984 = _RAND_1984[31:0];
  _RAND_1985 = {1{`RANDOM}};
  reg_csr_1985 = _RAND_1985[31:0];
  _RAND_1986 = {1{`RANDOM}};
  reg_csr_1986 = _RAND_1986[31:0];
  _RAND_1987 = {1{`RANDOM}};
  reg_csr_1987 = _RAND_1987[31:0];
  _RAND_1988 = {1{`RANDOM}};
  reg_csr_1988 = _RAND_1988[31:0];
  _RAND_1989 = {1{`RANDOM}};
  reg_csr_1989 = _RAND_1989[31:0];
  _RAND_1990 = {1{`RANDOM}};
  reg_csr_1990 = _RAND_1990[31:0];
  _RAND_1991 = {1{`RANDOM}};
  reg_csr_1991 = _RAND_1991[31:0];
  _RAND_1992 = {1{`RANDOM}};
  reg_csr_1992 = _RAND_1992[31:0];
  _RAND_1993 = {1{`RANDOM}};
  reg_csr_1993 = _RAND_1993[31:0];
  _RAND_1994 = {1{`RANDOM}};
  reg_csr_1994 = _RAND_1994[31:0];
  _RAND_1995 = {1{`RANDOM}};
  reg_csr_1995 = _RAND_1995[31:0];
  _RAND_1996 = {1{`RANDOM}};
  reg_csr_1996 = _RAND_1996[31:0];
  _RAND_1997 = {1{`RANDOM}};
  reg_csr_1997 = _RAND_1997[31:0];
  _RAND_1998 = {1{`RANDOM}};
  reg_csr_1998 = _RAND_1998[31:0];
  _RAND_1999 = {1{`RANDOM}};
  reg_csr_1999 = _RAND_1999[31:0];
  _RAND_2000 = {1{`RANDOM}};
  reg_csr_2000 = _RAND_2000[31:0];
  _RAND_2001 = {1{`RANDOM}};
  reg_csr_2001 = _RAND_2001[31:0];
  _RAND_2002 = {1{`RANDOM}};
  reg_csr_2002 = _RAND_2002[31:0];
  _RAND_2003 = {1{`RANDOM}};
  reg_csr_2003 = _RAND_2003[31:0];
  _RAND_2004 = {1{`RANDOM}};
  reg_csr_2004 = _RAND_2004[31:0];
  _RAND_2005 = {1{`RANDOM}};
  reg_csr_2005 = _RAND_2005[31:0];
  _RAND_2006 = {1{`RANDOM}};
  reg_csr_2006 = _RAND_2006[31:0];
  _RAND_2007 = {1{`RANDOM}};
  reg_csr_2007 = _RAND_2007[31:0];
  _RAND_2008 = {1{`RANDOM}};
  reg_csr_2008 = _RAND_2008[31:0];
  _RAND_2009 = {1{`RANDOM}};
  reg_csr_2009 = _RAND_2009[31:0];
  _RAND_2010 = {1{`RANDOM}};
  reg_csr_2010 = _RAND_2010[31:0];
  _RAND_2011 = {1{`RANDOM}};
  reg_csr_2011 = _RAND_2011[31:0];
  _RAND_2012 = {1{`RANDOM}};
  reg_csr_2012 = _RAND_2012[31:0];
  _RAND_2013 = {1{`RANDOM}};
  reg_csr_2013 = _RAND_2013[31:0];
  _RAND_2014 = {1{`RANDOM}};
  reg_csr_2014 = _RAND_2014[31:0];
  _RAND_2015 = {1{`RANDOM}};
  reg_csr_2015 = _RAND_2015[31:0];
  _RAND_2016 = {1{`RANDOM}};
  reg_csr_2016 = _RAND_2016[31:0];
  _RAND_2017 = {1{`RANDOM}};
  reg_csr_2017 = _RAND_2017[31:0];
  _RAND_2018 = {1{`RANDOM}};
  reg_csr_2018 = _RAND_2018[31:0];
  _RAND_2019 = {1{`RANDOM}};
  reg_csr_2019 = _RAND_2019[31:0];
  _RAND_2020 = {1{`RANDOM}};
  reg_csr_2020 = _RAND_2020[31:0];
  _RAND_2021 = {1{`RANDOM}};
  reg_csr_2021 = _RAND_2021[31:0];
  _RAND_2022 = {1{`RANDOM}};
  reg_csr_2022 = _RAND_2022[31:0];
  _RAND_2023 = {1{`RANDOM}};
  reg_csr_2023 = _RAND_2023[31:0];
  _RAND_2024 = {1{`RANDOM}};
  reg_csr_2024 = _RAND_2024[31:0];
  _RAND_2025 = {1{`RANDOM}};
  reg_csr_2025 = _RAND_2025[31:0];
  _RAND_2026 = {1{`RANDOM}};
  reg_csr_2026 = _RAND_2026[31:0];
  _RAND_2027 = {1{`RANDOM}};
  reg_csr_2027 = _RAND_2027[31:0];
  _RAND_2028 = {1{`RANDOM}};
  reg_csr_2028 = _RAND_2028[31:0];
  _RAND_2029 = {1{`RANDOM}};
  reg_csr_2029 = _RAND_2029[31:0];
  _RAND_2030 = {1{`RANDOM}};
  reg_csr_2030 = _RAND_2030[31:0];
  _RAND_2031 = {1{`RANDOM}};
  reg_csr_2031 = _RAND_2031[31:0];
  _RAND_2032 = {1{`RANDOM}};
  reg_csr_2032 = _RAND_2032[31:0];
  _RAND_2033 = {1{`RANDOM}};
  reg_csr_2033 = _RAND_2033[31:0];
  _RAND_2034 = {1{`RANDOM}};
  reg_csr_2034 = _RAND_2034[31:0];
  _RAND_2035 = {1{`RANDOM}};
  reg_csr_2035 = _RAND_2035[31:0];
  _RAND_2036 = {1{`RANDOM}};
  reg_csr_2036 = _RAND_2036[31:0];
  _RAND_2037 = {1{`RANDOM}};
  reg_csr_2037 = _RAND_2037[31:0];
  _RAND_2038 = {1{`RANDOM}};
  reg_csr_2038 = _RAND_2038[31:0];
  _RAND_2039 = {1{`RANDOM}};
  reg_csr_2039 = _RAND_2039[31:0];
  _RAND_2040 = {1{`RANDOM}};
  reg_csr_2040 = _RAND_2040[31:0];
  _RAND_2041 = {1{`RANDOM}};
  reg_csr_2041 = _RAND_2041[31:0];
  _RAND_2042 = {1{`RANDOM}};
  reg_csr_2042 = _RAND_2042[31:0];
  _RAND_2043 = {1{`RANDOM}};
  reg_csr_2043 = _RAND_2043[31:0];
  _RAND_2044 = {1{`RANDOM}};
  reg_csr_2044 = _RAND_2044[31:0];
  _RAND_2045 = {1{`RANDOM}};
  reg_csr_2045 = _RAND_2045[31:0];
  _RAND_2046 = {1{`RANDOM}};
  reg_csr_2046 = _RAND_2046[31:0];
  _RAND_2047 = {1{`RANDOM}};
  reg_csr_2047 = _RAND_2047[31:0];
  _RAND_2048 = {1{`RANDOM}};
  reg_csr_2048 = _RAND_2048[31:0];
  _RAND_2049 = {1{`RANDOM}};
  reg_csr_2049 = _RAND_2049[31:0];
  _RAND_2050 = {1{`RANDOM}};
  reg_csr_2050 = _RAND_2050[31:0];
  _RAND_2051 = {1{`RANDOM}};
  reg_csr_2051 = _RAND_2051[31:0];
  _RAND_2052 = {1{`RANDOM}};
  reg_csr_2052 = _RAND_2052[31:0];
  _RAND_2053 = {1{`RANDOM}};
  reg_csr_2053 = _RAND_2053[31:0];
  _RAND_2054 = {1{`RANDOM}};
  reg_csr_2054 = _RAND_2054[31:0];
  _RAND_2055 = {1{`RANDOM}};
  reg_csr_2055 = _RAND_2055[31:0];
  _RAND_2056 = {1{`RANDOM}};
  reg_csr_2056 = _RAND_2056[31:0];
  _RAND_2057 = {1{`RANDOM}};
  reg_csr_2057 = _RAND_2057[31:0];
  _RAND_2058 = {1{`RANDOM}};
  reg_csr_2058 = _RAND_2058[31:0];
  _RAND_2059 = {1{`RANDOM}};
  reg_csr_2059 = _RAND_2059[31:0];
  _RAND_2060 = {1{`RANDOM}};
  reg_csr_2060 = _RAND_2060[31:0];
  _RAND_2061 = {1{`RANDOM}};
  reg_csr_2061 = _RAND_2061[31:0];
  _RAND_2062 = {1{`RANDOM}};
  reg_csr_2062 = _RAND_2062[31:0];
  _RAND_2063 = {1{`RANDOM}};
  reg_csr_2063 = _RAND_2063[31:0];
  _RAND_2064 = {1{`RANDOM}};
  reg_csr_2064 = _RAND_2064[31:0];
  _RAND_2065 = {1{`RANDOM}};
  reg_csr_2065 = _RAND_2065[31:0];
  _RAND_2066 = {1{`RANDOM}};
  reg_csr_2066 = _RAND_2066[31:0];
  _RAND_2067 = {1{`RANDOM}};
  reg_csr_2067 = _RAND_2067[31:0];
  _RAND_2068 = {1{`RANDOM}};
  reg_csr_2068 = _RAND_2068[31:0];
  _RAND_2069 = {1{`RANDOM}};
  reg_csr_2069 = _RAND_2069[31:0];
  _RAND_2070 = {1{`RANDOM}};
  reg_csr_2070 = _RAND_2070[31:0];
  _RAND_2071 = {1{`RANDOM}};
  reg_csr_2071 = _RAND_2071[31:0];
  _RAND_2072 = {1{`RANDOM}};
  reg_csr_2072 = _RAND_2072[31:0];
  _RAND_2073 = {1{`RANDOM}};
  reg_csr_2073 = _RAND_2073[31:0];
  _RAND_2074 = {1{`RANDOM}};
  reg_csr_2074 = _RAND_2074[31:0];
  _RAND_2075 = {1{`RANDOM}};
  reg_csr_2075 = _RAND_2075[31:0];
  _RAND_2076 = {1{`RANDOM}};
  reg_csr_2076 = _RAND_2076[31:0];
  _RAND_2077 = {1{`RANDOM}};
  reg_csr_2077 = _RAND_2077[31:0];
  _RAND_2078 = {1{`RANDOM}};
  reg_csr_2078 = _RAND_2078[31:0];
  _RAND_2079 = {1{`RANDOM}};
  reg_csr_2079 = _RAND_2079[31:0];
  _RAND_2080 = {1{`RANDOM}};
  reg_csr_2080 = _RAND_2080[31:0];
  _RAND_2081 = {1{`RANDOM}};
  reg_csr_2081 = _RAND_2081[31:0];
  _RAND_2082 = {1{`RANDOM}};
  reg_csr_2082 = _RAND_2082[31:0];
  _RAND_2083 = {1{`RANDOM}};
  reg_csr_2083 = _RAND_2083[31:0];
  _RAND_2084 = {1{`RANDOM}};
  reg_csr_2084 = _RAND_2084[31:0];
  _RAND_2085 = {1{`RANDOM}};
  reg_csr_2085 = _RAND_2085[31:0];
  _RAND_2086 = {1{`RANDOM}};
  reg_csr_2086 = _RAND_2086[31:0];
  _RAND_2087 = {1{`RANDOM}};
  reg_csr_2087 = _RAND_2087[31:0];
  _RAND_2088 = {1{`RANDOM}};
  reg_csr_2088 = _RAND_2088[31:0];
  _RAND_2089 = {1{`RANDOM}};
  reg_csr_2089 = _RAND_2089[31:0];
  _RAND_2090 = {1{`RANDOM}};
  reg_csr_2090 = _RAND_2090[31:0];
  _RAND_2091 = {1{`RANDOM}};
  reg_csr_2091 = _RAND_2091[31:0];
  _RAND_2092 = {1{`RANDOM}};
  reg_csr_2092 = _RAND_2092[31:0];
  _RAND_2093 = {1{`RANDOM}};
  reg_csr_2093 = _RAND_2093[31:0];
  _RAND_2094 = {1{`RANDOM}};
  reg_csr_2094 = _RAND_2094[31:0];
  _RAND_2095 = {1{`RANDOM}};
  reg_csr_2095 = _RAND_2095[31:0];
  _RAND_2096 = {1{`RANDOM}};
  reg_csr_2096 = _RAND_2096[31:0];
  _RAND_2097 = {1{`RANDOM}};
  reg_csr_2097 = _RAND_2097[31:0];
  _RAND_2098 = {1{`RANDOM}};
  reg_csr_2098 = _RAND_2098[31:0];
  _RAND_2099 = {1{`RANDOM}};
  reg_csr_2099 = _RAND_2099[31:0];
  _RAND_2100 = {1{`RANDOM}};
  reg_csr_2100 = _RAND_2100[31:0];
  _RAND_2101 = {1{`RANDOM}};
  reg_csr_2101 = _RAND_2101[31:0];
  _RAND_2102 = {1{`RANDOM}};
  reg_csr_2102 = _RAND_2102[31:0];
  _RAND_2103 = {1{`RANDOM}};
  reg_csr_2103 = _RAND_2103[31:0];
  _RAND_2104 = {1{`RANDOM}};
  reg_csr_2104 = _RAND_2104[31:0];
  _RAND_2105 = {1{`RANDOM}};
  reg_csr_2105 = _RAND_2105[31:0];
  _RAND_2106 = {1{`RANDOM}};
  reg_csr_2106 = _RAND_2106[31:0];
  _RAND_2107 = {1{`RANDOM}};
  reg_csr_2107 = _RAND_2107[31:0];
  _RAND_2108 = {1{`RANDOM}};
  reg_csr_2108 = _RAND_2108[31:0];
  _RAND_2109 = {1{`RANDOM}};
  reg_csr_2109 = _RAND_2109[31:0];
  _RAND_2110 = {1{`RANDOM}};
  reg_csr_2110 = _RAND_2110[31:0];
  _RAND_2111 = {1{`RANDOM}};
  reg_csr_2111 = _RAND_2111[31:0];
  _RAND_2112 = {1{`RANDOM}};
  reg_csr_2112 = _RAND_2112[31:0];
  _RAND_2113 = {1{`RANDOM}};
  reg_csr_2113 = _RAND_2113[31:0];
  _RAND_2114 = {1{`RANDOM}};
  reg_csr_2114 = _RAND_2114[31:0];
  _RAND_2115 = {1{`RANDOM}};
  reg_csr_2115 = _RAND_2115[31:0];
  _RAND_2116 = {1{`RANDOM}};
  reg_csr_2116 = _RAND_2116[31:0];
  _RAND_2117 = {1{`RANDOM}};
  reg_csr_2117 = _RAND_2117[31:0];
  _RAND_2118 = {1{`RANDOM}};
  reg_csr_2118 = _RAND_2118[31:0];
  _RAND_2119 = {1{`RANDOM}};
  reg_csr_2119 = _RAND_2119[31:0];
  _RAND_2120 = {1{`RANDOM}};
  reg_csr_2120 = _RAND_2120[31:0];
  _RAND_2121 = {1{`RANDOM}};
  reg_csr_2121 = _RAND_2121[31:0];
  _RAND_2122 = {1{`RANDOM}};
  reg_csr_2122 = _RAND_2122[31:0];
  _RAND_2123 = {1{`RANDOM}};
  reg_csr_2123 = _RAND_2123[31:0];
  _RAND_2124 = {1{`RANDOM}};
  reg_csr_2124 = _RAND_2124[31:0];
  _RAND_2125 = {1{`RANDOM}};
  reg_csr_2125 = _RAND_2125[31:0];
  _RAND_2126 = {1{`RANDOM}};
  reg_csr_2126 = _RAND_2126[31:0];
  _RAND_2127 = {1{`RANDOM}};
  reg_csr_2127 = _RAND_2127[31:0];
  _RAND_2128 = {1{`RANDOM}};
  reg_csr_2128 = _RAND_2128[31:0];
  _RAND_2129 = {1{`RANDOM}};
  reg_csr_2129 = _RAND_2129[31:0];
  _RAND_2130 = {1{`RANDOM}};
  reg_csr_2130 = _RAND_2130[31:0];
  _RAND_2131 = {1{`RANDOM}};
  reg_csr_2131 = _RAND_2131[31:0];
  _RAND_2132 = {1{`RANDOM}};
  reg_csr_2132 = _RAND_2132[31:0];
  _RAND_2133 = {1{`RANDOM}};
  reg_csr_2133 = _RAND_2133[31:0];
  _RAND_2134 = {1{`RANDOM}};
  reg_csr_2134 = _RAND_2134[31:0];
  _RAND_2135 = {1{`RANDOM}};
  reg_csr_2135 = _RAND_2135[31:0];
  _RAND_2136 = {1{`RANDOM}};
  reg_csr_2136 = _RAND_2136[31:0];
  _RAND_2137 = {1{`RANDOM}};
  reg_csr_2137 = _RAND_2137[31:0];
  _RAND_2138 = {1{`RANDOM}};
  reg_csr_2138 = _RAND_2138[31:0];
  _RAND_2139 = {1{`RANDOM}};
  reg_csr_2139 = _RAND_2139[31:0];
  _RAND_2140 = {1{`RANDOM}};
  reg_csr_2140 = _RAND_2140[31:0];
  _RAND_2141 = {1{`RANDOM}};
  reg_csr_2141 = _RAND_2141[31:0];
  _RAND_2142 = {1{`RANDOM}};
  reg_csr_2142 = _RAND_2142[31:0];
  _RAND_2143 = {1{`RANDOM}};
  reg_csr_2143 = _RAND_2143[31:0];
  _RAND_2144 = {1{`RANDOM}};
  reg_csr_2144 = _RAND_2144[31:0];
  _RAND_2145 = {1{`RANDOM}};
  reg_csr_2145 = _RAND_2145[31:0];
  _RAND_2146 = {1{`RANDOM}};
  reg_csr_2146 = _RAND_2146[31:0];
  _RAND_2147 = {1{`RANDOM}};
  reg_csr_2147 = _RAND_2147[31:0];
  _RAND_2148 = {1{`RANDOM}};
  reg_csr_2148 = _RAND_2148[31:0];
  _RAND_2149 = {1{`RANDOM}};
  reg_csr_2149 = _RAND_2149[31:0];
  _RAND_2150 = {1{`RANDOM}};
  reg_csr_2150 = _RAND_2150[31:0];
  _RAND_2151 = {1{`RANDOM}};
  reg_csr_2151 = _RAND_2151[31:0];
  _RAND_2152 = {1{`RANDOM}};
  reg_csr_2152 = _RAND_2152[31:0];
  _RAND_2153 = {1{`RANDOM}};
  reg_csr_2153 = _RAND_2153[31:0];
  _RAND_2154 = {1{`RANDOM}};
  reg_csr_2154 = _RAND_2154[31:0];
  _RAND_2155 = {1{`RANDOM}};
  reg_csr_2155 = _RAND_2155[31:0];
  _RAND_2156 = {1{`RANDOM}};
  reg_csr_2156 = _RAND_2156[31:0];
  _RAND_2157 = {1{`RANDOM}};
  reg_csr_2157 = _RAND_2157[31:0];
  _RAND_2158 = {1{`RANDOM}};
  reg_csr_2158 = _RAND_2158[31:0];
  _RAND_2159 = {1{`RANDOM}};
  reg_csr_2159 = _RAND_2159[31:0];
  _RAND_2160 = {1{`RANDOM}};
  reg_csr_2160 = _RAND_2160[31:0];
  _RAND_2161 = {1{`RANDOM}};
  reg_csr_2161 = _RAND_2161[31:0];
  _RAND_2162 = {1{`RANDOM}};
  reg_csr_2162 = _RAND_2162[31:0];
  _RAND_2163 = {1{`RANDOM}};
  reg_csr_2163 = _RAND_2163[31:0];
  _RAND_2164 = {1{`RANDOM}};
  reg_csr_2164 = _RAND_2164[31:0];
  _RAND_2165 = {1{`RANDOM}};
  reg_csr_2165 = _RAND_2165[31:0];
  _RAND_2166 = {1{`RANDOM}};
  reg_csr_2166 = _RAND_2166[31:0];
  _RAND_2167 = {1{`RANDOM}};
  reg_csr_2167 = _RAND_2167[31:0];
  _RAND_2168 = {1{`RANDOM}};
  reg_csr_2168 = _RAND_2168[31:0];
  _RAND_2169 = {1{`RANDOM}};
  reg_csr_2169 = _RAND_2169[31:0];
  _RAND_2170 = {1{`RANDOM}};
  reg_csr_2170 = _RAND_2170[31:0];
  _RAND_2171 = {1{`RANDOM}};
  reg_csr_2171 = _RAND_2171[31:0];
  _RAND_2172 = {1{`RANDOM}};
  reg_csr_2172 = _RAND_2172[31:0];
  _RAND_2173 = {1{`RANDOM}};
  reg_csr_2173 = _RAND_2173[31:0];
  _RAND_2174 = {1{`RANDOM}};
  reg_csr_2174 = _RAND_2174[31:0];
  _RAND_2175 = {1{`RANDOM}};
  reg_csr_2175 = _RAND_2175[31:0];
  _RAND_2176 = {1{`RANDOM}};
  reg_csr_2176 = _RAND_2176[31:0];
  _RAND_2177 = {1{`RANDOM}};
  reg_csr_2177 = _RAND_2177[31:0];
  _RAND_2178 = {1{`RANDOM}};
  reg_csr_2178 = _RAND_2178[31:0];
  _RAND_2179 = {1{`RANDOM}};
  reg_csr_2179 = _RAND_2179[31:0];
  _RAND_2180 = {1{`RANDOM}};
  reg_csr_2180 = _RAND_2180[31:0];
  _RAND_2181 = {1{`RANDOM}};
  reg_csr_2181 = _RAND_2181[31:0];
  _RAND_2182 = {1{`RANDOM}};
  reg_csr_2182 = _RAND_2182[31:0];
  _RAND_2183 = {1{`RANDOM}};
  reg_csr_2183 = _RAND_2183[31:0];
  _RAND_2184 = {1{`RANDOM}};
  reg_csr_2184 = _RAND_2184[31:0];
  _RAND_2185 = {1{`RANDOM}};
  reg_csr_2185 = _RAND_2185[31:0];
  _RAND_2186 = {1{`RANDOM}};
  reg_csr_2186 = _RAND_2186[31:0];
  _RAND_2187 = {1{`RANDOM}};
  reg_csr_2187 = _RAND_2187[31:0];
  _RAND_2188 = {1{`RANDOM}};
  reg_csr_2188 = _RAND_2188[31:0];
  _RAND_2189 = {1{`RANDOM}};
  reg_csr_2189 = _RAND_2189[31:0];
  _RAND_2190 = {1{`RANDOM}};
  reg_csr_2190 = _RAND_2190[31:0];
  _RAND_2191 = {1{`RANDOM}};
  reg_csr_2191 = _RAND_2191[31:0];
  _RAND_2192 = {1{`RANDOM}};
  reg_csr_2192 = _RAND_2192[31:0];
  _RAND_2193 = {1{`RANDOM}};
  reg_csr_2193 = _RAND_2193[31:0];
  _RAND_2194 = {1{`RANDOM}};
  reg_csr_2194 = _RAND_2194[31:0];
  _RAND_2195 = {1{`RANDOM}};
  reg_csr_2195 = _RAND_2195[31:0];
  _RAND_2196 = {1{`RANDOM}};
  reg_csr_2196 = _RAND_2196[31:0];
  _RAND_2197 = {1{`RANDOM}};
  reg_csr_2197 = _RAND_2197[31:0];
  _RAND_2198 = {1{`RANDOM}};
  reg_csr_2198 = _RAND_2198[31:0];
  _RAND_2199 = {1{`RANDOM}};
  reg_csr_2199 = _RAND_2199[31:0];
  _RAND_2200 = {1{`RANDOM}};
  reg_csr_2200 = _RAND_2200[31:0];
  _RAND_2201 = {1{`RANDOM}};
  reg_csr_2201 = _RAND_2201[31:0];
  _RAND_2202 = {1{`RANDOM}};
  reg_csr_2202 = _RAND_2202[31:0];
  _RAND_2203 = {1{`RANDOM}};
  reg_csr_2203 = _RAND_2203[31:0];
  _RAND_2204 = {1{`RANDOM}};
  reg_csr_2204 = _RAND_2204[31:0];
  _RAND_2205 = {1{`RANDOM}};
  reg_csr_2205 = _RAND_2205[31:0];
  _RAND_2206 = {1{`RANDOM}};
  reg_csr_2206 = _RAND_2206[31:0];
  _RAND_2207 = {1{`RANDOM}};
  reg_csr_2207 = _RAND_2207[31:0];
  _RAND_2208 = {1{`RANDOM}};
  reg_csr_2208 = _RAND_2208[31:0];
  _RAND_2209 = {1{`RANDOM}};
  reg_csr_2209 = _RAND_2209[31:0];
  _RAND_2210 = {1{`RANDOM}};
  reg_csr_2210 = _RAND_2210[31:0];
  _RAND_2211 = {1{`RANDOM}};
  reg_csr_2211 = _RAND_2211[31:0];
  _RAND_2212 = {1{`RANDOM}};
  reg_csr_2212 = _RAND_2212[31:0];
  _RAND_2213 = {1{`RANDOM}};
  reg_csr_2213 = _RAND_2213[31:0];
  _RAND_2214 = {1{`RANDOM}};
  reg_csr_2214 = _RAND_2214[31:0];
  _RAND_2215 = {1{`RANDOM}};
  reg_csr_2215 = _RAND_2215[31:0];
  _RAND_2216 = {1{`RANDOM}};
  reg_csr_2216 = _RAND_2216[31:0];
  _RAND_2217 = {1{`RANDOM}};
  reg_csr_2217 = _RAND_2217[31:0];
  _RAND_2218 = {1{`RANDOM}};
  reg_csr_2218 = _RAND_2218[31:0];
  _RAND_2219 = {1{`RANDOM}};
  reg_csr_2219 = _RAND_2219[31:0];
  _RAND_2220 = {1{`RANDOM}};
  reg_csr_2220 = _RAND_2220[31:0];
  _RAND_2221 = {1{`RANDOM}};
  reg_csr_2221 = _RAND_2221[31:0];
  _RAND_2222 = {1{`RANDOM}};
  reg_csr_2222 = _RAND_2222[31:0];
  _RAND_2223 = {1{`RANDOM}};
  reg_csr_2223 = _RAND_2223[31:0];
  _RAND_2224 = {1{`RANDOM}};
  reg_csr_2224 = _RAND_2224[31:0];
  _RAND_2225 = {1{`RANDOM}};
  reg_csr_2225 = _RAND_2225[31:0];
  _RAND_2226 = {1{`RANDOM}};
  reg_csr_2226 = _RAND_2226[31:0];
  _RAND_2227 = {1{`RANDOM}};
  reg_csr_2227 = _RAND_2227[31:0];
  _RAND_2228 = {1{`RANDOM}};
  reg_csr_2228 = _RAND_2228[31:0];
  _RAND_2229 = {1{`RANDOM}};
  reg_csr_2229 = _RAND_2229[31:0];
  _RAND_2230 = {1{`RANDOM}};
  reg_csr_2230 = _RAND_2230[31:0];
  _RAND_2231 = {1{`RANDOM}};
  reg_csr_2231 = _RAND_2231[31:0];
  _RAND_2232 = {1{`RANDOM}};
  reg_csr_2232 = _RAND_2232[31:0];
  _RAND_2233 = {1{`RANDOM}};
  reg_csr_2233 = _RAND_2233[31:0];
  _RAND_2234 = {1{`RANDOM}};
  reg_csr_2234 = _RAND_2234[31:0];
  _RAND_2235 = {1{`RANDOM}};
  reg_csr_2235 = _RAND_2235[31:0];
  _RAND_2236 = {1{`RANDOM}};
  reg_csr_2236 = _RAND_2236[31:0];
  _RAND_2237 = {1{`RANDOM}};
  reg_csr_2237 = _RAND_2237[31:0];
  _RAND_2238 = {1{`RANDOM}};
  reg_csr_2238 = _RAND_2238[31:0];
  _RAND_2239 = {1{`RANDOM}};
  reg_csr_2239 = _RAND_2239[31:0];
  _RAND_2240 = {1{`RANDOM}};
  reg_csr_2240 = _RAND_2240[31:0];
  _RAND_2241 = {1{`RANDOM}};
  reg_csr_2241 = _RAND_2241[31:0];
  _RAND_2242 = {1{`RANDOM}};
  reg_csr_2242 = _RAND_2242[31:0];
  _RAND_2243 = {1{`RANDOM}};
  reg_csr_2243 = _RAND_2243[31:0];
  _RAND_2244 = {1{`RANDOM}};
  reg_csr_2244 = _RAND_2244[31:0];
  _RAND_2245 = {1{`RANDOM}};
  reg_csr_2245 = _RAND_2245[31:0];
  _RAND_2246 = {1{`RANDOM}};
  reg_csr_2246 = _RAND_2246[31:0];
  _RAND_2247 = {1{`RANDOM}};
  reg_csr_2247 = _RAND_2247[31:0];
  _RAND_2248 = {1{`RANDOM}};
  reg_csr_2248 = _RAND_2248[31:0];
  _RAND_2249 = {1{`RANDOM}};
  reg_csr_2249 = _RAND_2249[31:0];
  _RAND_2250 = {1{`RANDOM}};
  reg_csr_2250 = _RAND_2250[31:0];
  _RAND_2251 = {1{`RANDOM}};
  reg_csr_2251 = _RAND_2251[31:0];
  _RAND_2252 = {1{`RANDOM}};
  reg_csr_2252 = _RAND_2252[31:0];
  _RAND_2253 = {1{`RANDOM}};
  reg_csr_2253 = _RAND_2253[31:0];
  _RAND_2254 = {1{`RANDOM}};
  reg_csr_2254 = _RAND_2254[31:0];
  _RAND_2255 = {1{`RANDOM}};
  reg_csr_2255 = _RAND_2255[31:0];
  _RAND_2256 = {1{`RANDOM}};
  reg_csr_2256 = _RAND_2256[31:0];
  _RAND_2257 = {1{`RANDOM}};
  reg_csr_2257 = _RAND_2257[31:0];
  _RAND_2258 = {1{`RANDOM}};
  reg_csr_2258 = _RAND_2258[31:0];
  _RAND_2259 = {1{`RANDOM}};
  reg_csr_2259 = _RAND_2259[31:0];
  _RAND_2260 = {1{`RANDOM}};
  reg_csr_2260 = _RAND_2260[31:0];
  _RAND_2261 = {1{`RANDOM}};
  reg_csr_2261 = _RAND_2261[31:0];
  _RAND_2262 = {1{`RANDOM}};
  reg_csr_2262 = _RAND_2262[31:0];
  _RAND_2263 = {1{`RANDOM}};
  reg_csr_2263 = _RAND_2263[31:0];
  _RAND_2264 = {1{`RANDOM}};
  reg_csr_2264 = _RAND_2264[31:0];
  _RAND_2265 = {1{`RANDOM}};
  reg_csr_2265 = _RAND_2265[31:0];
  _RAND_2266 = {1{`RANDOM}};
  reg_csr_2266 = _RAND_2266[31:0];
  _RAND_2267 = {1{`RANDOM}};
  reg_csr_2267 = _RAND_2267[31:0];
  _RAND_2268 = {1{`RANDOM}};
  reg_csr_2268 = _RAND_2268[31:0];
  _RAND_2269 = {1{`RANDOM}};
  reg_csr_2269 = _RAND_2269[31:0];
  _RAND_2270 = {1{`RANDOM}};
  reg_csr_2270 = _RAND_2270[31:0];
  _RAND_2271 = {1{`RANDOM}};
  reg_csr_2271 = _RAND_2271[31:0];
  _RAND_2272 = {1{`RANDOM}};
  reg_csr_2272 = _RAND_2272[31:0];
  _RAND_2273 = {1{`RANDOM}};
  reg_csr_2273 = _RAND_2273[31:0];
  _RAND_2274 = {1{`RANDOM}};
  reg_csr_2274 = _RAND_2274[31:0];
  _RAND_2275 = {1{`RANDOM}};
  reg_csr_2275 = _RAND_2275[31:0];
  _RAND_2276 = {1{`RANDOM}};
  reg_csr_2276 = _RAND_2276[31:0];
  _RAND_2277 = {1{`RANDOM}};
  reg_csr_2277 = _RAND_2277[31:0];
  _RAND_2278 = {1{`RANDOM}};
  reg_csr_2278 = _RAND_2278[31:0];
  _RAND_2279 = {1{`RANDOM}};
  reg_csr_2279 = _RAND_2279[31:0];
  _RAND_2280 = {1{`RANDOM}};
  reg_csr_2280 = _RAND_2280[31:0];
  _RAND_2281 = {1{`RANDOM}};
  reg_csr_2281 = _RAND_2281[31:0];
  _RAND_2282 = {1{`RANDOM}};
  reg_csr_2282 = _RAND_2282[31:0];
  _RAND_2283 = {1{`RANDOM}};
  reg_csr_2283 = _RAND_2283[31:0];
  _RAND_2284 = {1{`RANDOM}};
  reg_csr_2284 = _RAND_2284[31:0];
  _RAND_2285 = {1{`RANDOM}};
  reg_csr_2285 = _RAND_2285[31:0];
  _RAND_2286 = {1{`RANDOM}};
  reg_csr_2286 = _RAND_2286[31:0];
  _RAND_2287 = {1{`RANDOM}};
  reg_csr_2287 = _RAND_2287[31:0];
  _RAND_2288 = {1{`RANDOM}};
  reg_csr_2288 = _RAND_2288[31:0];
  _RAND_2289 = {1{`RANDOM}};
  reg_csr_2289 = _RAND_2289[31:0];
  _RAND_2290 = {1{`RANDOM}};
  reg_csr_2290 = _RAND_2290[31:0];
  _RAND_2291 = {1{`RANDOM}};
  reg_csr_2291 = _RAND_2291[31:0];
  _RAND_2292 = {1{`RANDOM}};
  reg_csr_2292 = _RAND_2292[31:0];
  _RAND_2293 = {1{`RANDOM}};
  reg_csr_2293 = _RAND_2293[31:0];
  _RAND_2294 = {1{`RANDOM}};
  reg_csr_2294 = _RAND_2294[31:0];
  _RAND_2295 = {1{`RANDOM}};
  reg_csr_2295 = _RAND_2295[31:0];
  _RAND_2296 = {1{`RANDOM}};
  reg_csr_2296 = _RAND_2296[31:0];
  _RAND_2297 = {1{`RANDOM}};
  reg_csr_2297 = _RAND_2297[31:0];
  _RAND_2298 = {1{`RANDOM}};
  reg_csr_2298 = _RAND_2298[31:0];
  _RAND_2299 = {1{`RANDOM}};
  reg_csr_2299 = _RAND_2299[31:0];
  _RAND_2300 = {1{`RANDOM}};
  reg_csr_2300 = _RAND_2300[31:0];
  _RAND_2301 = {1{`RANDOM}};
  reg_csr_2301 = _RAND_2301[31:0];
  _RAND_2302 = {1{`RANDOM}};
  reg_csr_2302 = _RAND_2302[31:0];
  _RAND_2303 = {1{`RANDOM}};
  reg_csr_2303 = _RAND_2303[31:0];
  _RAND_2304 = {1{`RANDOM}};
  reg_csr_2304 = _RAND_2304[31:0];
  _RAND_2305 = {1{`RANDOM}};
  reg_csr_2305 = _RAND_2305[31:0];
  _RAND_2306 = {1{`RANDOM}};
  reg_csr_2306 = _RAND_2306[31:0];
  _RAND_2307 = {1{`RANDOM}};
  reg_csr_2307 = _RAND_2307[31:0];
  _RAND_2308 = {1{`RANDOM}};
  reg_csr_2308 = _RAND_2308[31:0];
  _RAND_2309 = {1{`RANDOM}};
  reg_csr_2309 = _RAND_2309[31:0];
  _RAND_2310 = {1{`RANDOM}};
  reg_csr_2310 = _RAND_2310[31:0];
  _RAND_2311 = {1{`RANDOM}};
  reg_csr_2311 = _RAND_2311[31:0];
  _RAND_2312 = {1{`RANDOM}};
  reg_csr_2312 = _RAND_2312[31:0];
  _RAND_2313 = {1{`RANDOM}};
  reg_csr_2313 = _RAND_2313[31:0];
  _RAND_2314 = {1{`RANDOM}};
  reg_csr_2314 = _RAND_2314[31:0];
  _RAND_2315 = {1{`RANDOM}};
  reg_csr_2315 = _RAND_2315[31:0];
  _RAND_2316 = {1{`RANDOM}};
  reg_csr_2316 = _RAND_2316[31:0];
  _RAND_2317 = {1{`RANDOM}};
  reg_csr_2317 = _RAND_2317[31:0];
  _RAND_2318 = {1{`RANDOM}};
  reg_csr_2318 = _RAND_2318[31:0];
  _RAND_2319 = {1{`RANDOM}};
  reg_csr_2319 = _RAND_2319[31:0];
  _RAND_2320 = {1{`RANDOM}};
  reg_csr_2320 = _RAND_2320[31:0];
  _RAND_2321 = {1{`RANDOM}};
  reg_csr_2321 = _RAND_2321[31:0];
  _RAND_2322 = {1{`RANDOM}};
  reg_csr_2322 = _RAND_2322[31:0];
  _RAND_2323 = {1{`RANDOM}};
  reg_csr_2323 = _RAND_2323[31:0];
  _RAND_2324 = {1{`RANDOM}};
  reg_csr_2324 = _RAND_2324[31:0];
  _RAND_2325 = {1{`RANDOM}};
  reg_csr_2325 = _RAND_2325[31:0];
  _RAND_2326 = {1{`RANDOM}};
  reg_csr_2326 = _RAND_2326[31:0];
  _RAND_2327 = {1{`RANDOM}};
  reg_csr_2327 = _RAND_2327[31:0];
  _RAND_2328 = {1{`RANDOM}};
  reg_csr_2328 = _RAND_2328[31:0];
  _RAND_2329 = {1{`RANDOM}};
  reg_csr_2329 = _RAND_2329[31:0];
  _RAND_2330 = {1{`RANDOM}};
  reg_csr_2330 = _RAND_2330[31:0];
  _RAND_2331 = {1{`RANDOM}};
  reg_csr_2331 = _RAND_2331[31:0];
  _RAND_2332 = {1{`RANDOM}};
  reg_csr_2332 = _RAND_2332[31:0];
  _RAND_2333 = {1{`RANDOM}};
  reg_csr_2333 = _RAND_2333[31:0];
  _RAND_2334 = {1{`RANDOM}};
  reg_csr_2334 = _RAND_2334[31:0];
  _RAND_2335 = {1{`RANDOM}};
  reg_csr_2335 = _RAND_2335[31:0];
  _RAND_2336 = {1{`RANDOM}};
  reg_csr_2336 = _RAND_2336[31:0];
  _RAND_2337 = {1{`RANDOM}};
  reg_csr_2337 = _RAND_2337[31:0];
  _RAND_2338 = {1{`RANDOM}};
  reg_csr_2338 = _RAND_2338[31:0];
  _RAND_2339 = {1{`RANDOM}};
  reg_csr_2339 = _RAND_2339[31:0];
  _RAND_2340 = {1{`RANDOM}};
  reg_csr_2340 = _RAND_2340[31:0];
  _RAND_2341 = {1{`RANDOM}};
  reg_csr_2341 = _RAND_2341[31:0];
  _RAND_2342 = {1{`RANDOM}};
  reg_csr_2342 = _RAND_2342[31:0];
  _RAND_2343 = {1{`RANDOM}};
  reg_csr_2343 = _RAND_2343[31:0];
  _RAND_2344 = {1{`RANDOM}};
  reg_csr_2344 = _RAND_2344[31:0];
  _RAND_2345 = {1{`RANDOM}};
  reg_csr_2345 = _RAND_2345[31:0];
  _RAND_2346 = {1{`RANDOM}};
  reg_csr_2346 = _RAND_2346[31:0];
  _RAND_2347 = {1{`RANDOM}};
  reg_csr_2347 = _RAND_2347[31:0];
  _RAND_2348 = {1{`RANDOM}};
  reg_csr_2348 = _RAND_2348[31:0];
  _RAND_2349 = {1{`RANDOM}};
  reg_csr_2349 = _RAND_2349[31:0];
  _RAND_2350 = {1{`RANDOM}};
  reg_csr_2350 = _RAND_2350[31:0];
  _RAND_2351 = {1{`RANDOM}};
  reg_csr_2351 = _RAND_2351[31:0];
  _RAND_2352 = {1{`RANDOM}};
  reg_csr_2352 = _RAND_2352[31:0];
  _RAND_2353 = {1{`RANDOM}};
  reg_csr_2353 = _RAND_2353[31:0];
  _RAND_2354 = {1{`RANDOM}};
  reg_csr_2354 = _RAND_2354[31:0];
  _RAND_2355 = {1{`RANDOM}};
  reg_csr_2355 = _RAND_2355[31:0];
  _RAND_2356 = {1{`RANDOM}};
  reg_csr_2356 = _RAND_2356[31:0];
  _RAND_2357 = {1{`RANDOM}};
  reg_csr_2357 = _RAND_2357[31:0];
  _RAND_2358 = {1{`RANDOM}};
  reg_csr_2358 = _RAND_2358[31:0];
  _RAND_2359 = {1{`RANDOM}};
  reg_csr_2359 = _RAND_2359[31:0];
  _RAND_2360 = {1{`RANDOM}};
  reg_csr_2360 = _RAND_2360[31:0];
  _RAND_2361 = {1{`RANDOM}};
  reg_csr_2361 = _RAND_2361[31:0];
  _RAND_2362 = {1{`RANDOM}};
  reg_csr_2362 = _RAND_2362[31:0];
  _RAND_2363 = {1{`RANDOM}};
  reg_csr_2363 = _RAND_2363[31:0];
  _RAND_2364 = {1{`RANDOM}};
  reg_csr_2364 = _RAND_2364[31:0];
  _RAND_2365 = {1{`RANDOM}};
  reg_csr_2365 = _RAND_2365[31:0];
  _RAND_2366 = {1{`RANDOM}};
  reg_csr_2366 = _RAND_2366[31:0];
  _RAND_2367 = {1{`RANDOM}};
  reg_csr_2367 = _RAND_2367[31:0];
  _RAND_2368 = {1{`RANDOM}};
  reg_csr_2368 = _RAND_2368[31:0];
  _RAND_2369 = {1{`RANDOM}};
  reg_csr_2369 = _RAND_2369[31:0];
  _RAND_2370 = {1{`RANDOM}};
  reg_csr_2370 = _RAND_2370[31:0];
  _RAND_2371 = {1{`RANDOM}};
  reg_csr_2371 = _RAND_2371[31:0];
  _RAND_2372 = {1{`RANDOM}};
  reg_csr_2372 = _RAND_2372[31:0];
  _RAND_2373 = {1{`RANDOM}};
  reg_csr_2373 = _RAND_2373[31:0];
  _RAND_2374 = {1{`RANDOM}};
  reg_csr_2374 = _RAND_2374[31:0];
  _RAND_2375 = {1{`RANDOM}};
  reg_csr_2375 = _RAND_2375[31:0];
  _RAND_2376 = {1{`RANDOM}};
  reg_csr_2376 = _RAND_2376[31:0];
  _RAND_2377 = {1{`RANDOM}};
  reg_csr_2377 = _RAND_2377[31:0];
  _RAND_2378 = {1{`RANDOM}};
  reg_csr_2378 = _RAND_2378[31:0];
  _RAND_2379 = {1{`RANDOM}};
  reg_csr_2379 = _RAND_2379[31:0];
  _RAND_2380 = {1{`RANDOM}};
  reg_csr_2380 = _RAND_2380[31:0];
  _RAND_2381 = {1{`RANDOM}};
  reg_csr_2381 = _RAND_2381[31:0];
  _RAND_2382 = {1{`RANDOM}};
  reg_csr_2382 = _RAND_2382[31:0];
  _RAND_2383 = {1{`RANDOM}};
  reg_csr_2383 = _RAND_2383[31:0];
  _RAND_2384 = {1{`RANDOM}};
  reg_csr_2384 = _RAND_2384[31:0];
  _RAND_2385 = {1{`RANDOM}};
  reg_csr_2385 = _RAND_2385[31:0];
  _RAND_2386 = {1{`RANDOM}};
  reg_csr_2386 = _RAND_2386[31:0];
  _RAND_2387 = {1{`RANDOM}};
  reg_csr_2387 = _RAND_2387[31:0];
  _RAND_2388 = {1{`RANDOM}};
  reg_csr_2388 = _RAND_2388[31:0];
  _RAND_2389 = {1{`RANDOM}};
  reg_csr_2389 = _RAND_2389[31:0];
  _RAND_2390 = {1{`RANDOM}};
  reg_csr_2390 = _RAND_2390[31:0];
  _RAND_2391 = {1{`RANDOM}};
  reg_csr_2391 = _RAND_2391[31:0];
  _RAND_2392 = {1{`RANDOM}};
  reg_csr_2392 = _RAND_2392[31:0];
  _RAND_2393 = {1{`RANDOM}};
  reg_csr_2393 = _RAND_2393[31:0];
  _RAND_2394 = {1{`RANDOM}};
  reg_csr_2394 = _RAND_2394[31:0];
  _RAND_2395 = {1{`RANDOM}};
  reg_csr_2395 = _RAND_2395[31:0];
  _RAND_2396 = {1{`RANDOM}};
  reg_csr_2396 = _RAND_2396[31:0];
  _RAND_2397 = {1{`RANDOM}};
  reg_csr_2397 = _RAND_2397[31:0];
  _RAND_2398 = {1{`RANDOM}};
  reg_csr_2398 = _RAND_2398[31:0];
  _RAND_2399 = {1{`RANDOM}};
  reg_csr_2399 = _RAND_2399[31:0];
  _RAND_2400 = {1{`RANDOM}};
  reg_csr_2400 = _RAND_2400[31:0];
  _RAND_2401 = {1{`RANDOM}};
  reg_csr_2401 = _RAND_2401[31:0];
  _RAND_2402 = {1{`RANDOM}};
  reg_csr_2402 = _RAND_2402[31:0];
  _RAND_2403 = {1{`RANDOM}};
  reg_csr_2403 = _RAND_2403[31:0];
  _RAND_2404 = {1{`RANDOM}};
  reg_csr_2404 = _RAND_2404[31:0];
  _RAND_2405 = {1{`RANDOM}};
  reg_csr_2405 = _RAND_2405[31:0];
  _RAND_2406 = {1{`RANDOM}};
  reg_csr_2406 = _RAND_2406[31:0];
  _RAND_2407 = {1{`RANDOM}};
  reg_csr_2407 = _RAND_2407[31:0];
  _RAND_2408 = {1{`RANDOM}};
  reg_csr_2408 = _RAND_2408[31:0];
  _RAND_2409 = {1{`RANDOM}};
  reg_csr_2409 = _RAND_2409[31:0];
  _RAND_2410 = {1{`RANDOM}};
  reg_csr_2410 = _RAND_2410[31:0];
  _RAND_2411 = {1{`RANDOM}};
  reg_csr_2411 = _RAND_2411[31:0];
  _RAND_2412 = {1{`RANDOM}};
  reg_csr_2412 = _RAND_2412[31:0];
  _RAND_2413 = {1{`RANDOM}};
  reg_csr_2413 = _RAND_2413[31:0];
  _RAND_2414 = {1{`RANDOM}};
  reg_csr_2414 = _RAND_2414[31:0];
  _RAND_2415 = {1{`RANDOM}};
  reg_csr_2415 = _RAND_2415[31:0];
  _RAND_2416 = {1{`RANDOM}};
  reg_csr_2416 = _RAND_2416[31:0];
  _RAND_2417 = {1{`RANDOM}};
  reg_csr_2417 = _RAND_2417[31:0];
  _RAND_2418 = {1{`RANDOM}};
  reg_csr_2418 = _RAND_2418[31:0];
  _RAND_2419 = {1{`RANDOM}};
  reg_csr_2419 = _RAND_2419[31:0];
  _RAND_2420 = {1{`RANDOM}};
  reg_csr_2420 = _RAND_2420[31:0];
  _RAND_2421 = {1{`RANDOM}};
  reg_csr_2421 = _RAND_2421[31:0];
  _RAND_2422 = {1{`RANDOM}};
  reg_csr_2422 = _RAND_2422[31:0];
  _RAND_2423 = {1{`RANDOM}};
  reg_csr_2423 = _RAND_2423[31:0];
  _RAND_2424 = {1{`RANDOM}};
  reg_csr_2424 = _RAND_2424[31:0];
  _RAND_2425 = {1{`RANDOM}};
  reg_csr_2425 = _RAND_2425[31:0];
  _RAND_2426 = {1{`RANDOM}};
  reg_csr_2426 = _RAND_2426[31:0];
  _RAND_2427 = {1{`RANDOM}};
  reg_csr_2427 = _RAND_2427[31:0];
  _RAND_2428 = {1{`RANDOM}};
  reg_csr_2428 = _RAND_2428[31:0];
  _RAND_2429 = {1{`RANDOM}};
  reg_csr_2429 = _RAND_2429[31:0];
  _RAND_2430 = {1{`RANDOM}};
  reg_csr_2430 = _RAND_2430[31:0];
  _RAND_2431 = {1{`RANDOM}};
  reg_csr_2431 = _RAND_2431[31:0];
  _RAND_2432 = {1{`RANDOM}};
  reg_csr_2432 = _RAND_2432[31:0];
  _RAND_2433 = {1{`RANDOM}};
  reg_csr_2433 = _RAND_2433[31:0];
  _RAND_2434 = {1{`RANDOM}};
  reg_csr_2434 = _RAND_2434[31:0];
  _RAND_2435 = {1{`RANDOM}};
  reg_csr_2435 = _RAND_2435[31:0];
  _RAND_2436 = {1{`RANDOM}};
  reg_csr_2436 = _RAND_2436[31:0];
  _RAND_2437 = {1{`RANDOM}};
  reg_csr_2437 = _RAND_2437[31:0];
  _RAND_2438 = {1{`RANDOM}};
  reg_csr_2438 = _RAND_2438[31:0];
  _RAND_2439 = {1{`RANDOM}};
  reg_csr_2439 = _RAND_2439[31:0];
  _RAND_2440 = {1{`RANDOM}};
  reg_csr_2440 = _RAND_2440[31:0];
  _RAND_2441 = {1{`RANDOM}};
  reg_csr_2441 = _RAND_2441[31:0];
  _RAND_2442 = {1{`RANDOM}};
  reg_csr_2442 = _RAND_2442[31:0];
  _RAND_2443 = {1{`RANDOM}};
  reg_csr_2443 = _RAND_2443[31:0];
  _RAND_2444 = {1{`RANDOM}};
  reg_csr_2444 = _RAND_2444[31:0];
  _RAND_2445 = {1{`RANDOM}};
  reg_csr_2445 = _RAND_2445[31:0];
  _RAND_2446 = {1{`RANDOM}};
  reg_csr_2446 = _RAND_2446[31:0];
  _RAND_2447 = {1{`RANDOM}};
  reg_csr_2447 = _RAND_2447[31:0];
  _RAND_2448 = {1{`RANDOM}};
  reg_csr_2448 = _RAND_2448[31:0];
  _RAND_2449 = {1{`RANDOM}};
  reg_csr_2449 = _RAND_2449[31:0];
  _RAND_2450 = {1{`RANDOM}};
  reg_csr_2450 = _RAND_2450[31:0];
  _RAND_2451 = {1{`RANDOM}};
  reg_csr_2451 = _RAND_2451[31:0];
  _RAND_2452 = {1{`RANDOM}};
  reg_csr_2452 = _RAND_2452[31:0];
  _RAND_2453 = {1{`RANDOM}};
  reg_csr_2453 = _RAND_2453[31:0];
  _RAND_2454 = {1{`RANDOM}};
  reg_csr_2454 = _RAND_2454[31:0];
  _RAND_2455 = {1{`RANDOM}};
  reg_csr_2455 = _RAND_2455[31:0];
  _RAND_2456 = {1{`RANDOM}};
  reg_csr_2456 = _RAND_2456[31:0];
  _RAND_2457 = {1{`RANDOM}};
  reg_csr_2457 = _RAND_2457[31:0];
  _RAND_2458 = {1{`RANDOM}};
  reg_csr_2458 = _RAND_2458[31:0];
  _RAND_2459 = {1{`RANDOM}};
  reg_csr_2459 = _RAND_2459[31:0];
  _RAND_2460 = {1{`RANDOM}};
  reg_csr_2460 = _RAND_2460[31:0];
  _RAND_2461 = {1{`RANDOM}};
  reg_csr_2461 = _RAND_2461[31:0];
  _RAND_2462 = {1{`RANDOM}};
  reg_csr_2462 = _RAND_2462[31:0];
  _RAND_2463 = {1{`RANDOM}};
  reg_csr_2463 = _RAND_2463[31:0];
  _RAND_2464 = {1{`RANDOM}};
  reg_csr_2464 = _RAND_2464[31:0];
  _RAND_2465 = {1{`RANDOM}};
  reg_csr_2465 = _RAND_2465[31:0];
  _RAND_2466 = {1{`RANDOM}};
  reg_csr_2466 = _RAND_2466[31:0];
  _RAND_2467 = {1{`RANDOM}};
  reg_csr_2467 = _RAND_2467[31:0];
  _RAND_2468 = {1{`RANDOM}};
  reg_csr_2468 = _RAND_2468[31:0];
  _RAND_2469 = {1{`RANDOM}};
  reg_csr_2469 = _RAND_2469[31:0];
  _RAND_2470 = {1{`RANDOM}};
  reg_csr_2470 = _RAND_2470[31:0];
  _RAND_2471 = {1{`RANDOM}};
  reg_csr_2471 = _RAND_2471[31:0];
  _RAND_2472 = {1{`RANDOM}};
  reg_csr_2472 = _RAND_2472[31:0];
  _RAND_2473 = {1{`RANDOM}};
  reg_csr_2473 = _RAND_2473[31:0];
  _RAND_2474 = {1{`RANDOM}};
  reg_csr_2474 = _RAND_2474[31:0];
  _RAND_2475 = {1{`RANDOM}};
  reg_csr_2475 = _RAND_2475[31:0];
  _RAND_2476 = {1{`RANDOM}};
  reg_csr_2476 = _RAND_2476[31:0];
  _RAND_2477 = {1{`RANDOM}};
  reg_csr_2477 = _RAND_2477[31:0];
  _RAND_2478 = {1{`RANDOM}};
  reg_csr_2478 = _RAND_2478[31:0];
  _RAND_2479 = {1{`RANDOM}};
  reg_csr_2479 = _RAND_2479[31:0];
  _RAND_2480 = {1{`RANDOM}};
  reg_csr_2480 = _RAND_2480[31:0];
  _RAND_2481 = {1{`RANDOM}};
  reg_csr_2481 = _RAND_2481[31:0];
  _RAND_2482 = {1{`RANDOM}};
  reg_csr_2482 = _RAND_2482[31:0];
  _RAND_2483 = {1{`RANDOM}};
  reg_csr_2483 = _RAND_2483[31:0];
  _RAND_2484 = {1{`RANDOM}};
  reg_csr_2484 = _RAND_2484[31:0];
  _RAND_2485 = {1{`RANDOM}};
  reg_csr_2485 = _RAND_2485[31:0];
  _RAND_2486 = {1{`RANDOM}};
  reg_csr_2486 = _RAND_2486[31:0];
  _RAND_2487 = {1{`RANDOM}};
  reg_csr_2487 = _RAND_2487[31:0];
  _RAND_2488 = {1{`RANDOM}};
  reg_csr_2488 = _RAND_2488[31:0];
  _RAND_2489 = {1{`RANDOM}};
  reg_csr_2489 = _RAND_2489[31:0];
  _RAND_2490 = {1{`RANDOM}};
  reg_csr_2490 = _RAND_2490[31:0];
  _RAND_2491 = {1{`RANDOM}};
  reg_csr_2491 = _RAND_2491[31:0];
  _RAND_2492 = {1{`RANDOM}};
  reg_csr_2492 = _RAND_2492[31:0];
  _RAND_2493 = {1{`RANDOM}};
  reg_csr_2493 = _RAND_2493[31:0];
  _RAND_2494 = {1{`RANDOM}};
  reg_csr_2494 = _RAND_2494[31:0];
  _RAND_2495 = {1{`RANDOM}};
  reg_csr_2495 = _RAND_2495[31:0];
  _RAND_2496 = {1{`RANDOM}};
  reg_csr_2496 = _RAND_2496[31:0];
  _RAND_2497 = {1{`RANDOM}};
  reg_csr_2497 = _RAND_2497[31:0];
  _RAND_2498 = {1{`RANDOM}};
  reg_csr_2498 = _RAND_2498[31:0];
  _RAND_2499 = {1{`RANDOM}};
  reg_csr_2499 = _RAND_2499[31:0];
  _RAND_2500 = {1{`RANDOM}};
  reg_csr_2500 = _RAND_2500[31:0];
  _RAND_2501 = {1{`RANDOM}};
  reg_csr_2501 = _RAND_2501[31:0];
  _RAND_2502 = {1{`RANDOM}};
  reg_csr_2502 = _RAND_2502[31:0];
  _RAND_2503 = {1{`RANDOM}};
  reg_csr_2503 = _RAND_2503[31:0];
  _RAND_2504 = {1{`RANDOM}};
  reg_csr_2504 = _RAND_2504[31:0];
  _RAND_2505 = {1{`RANDOM}};
  reg_csr_2505 = _RAND_2505[31:0];
  _RAND_2506 = {1{`RANDOM}};
  reg_csr_2506 = _RAND_2506[31:0];
  _RAND_2507 = {1{`RANDOM}};
  reg_csr_2507 = _RAND_2507[31:0];
  _RAND_2508 = {1{`RANDOM}};
  reg_csr_2508 = _RAND_2508[31:0];
  _RAND_2509 = {1{`RANDOM}};
  reg_csr_2509 = _RAND_2509[31:0];
  _RAND_2510 = {1{`RANDOM}};
  reg_csr_2510 = _RAND_2510[31:0];
  _RAND_2511 = {1{`RANDOM}};
  reg_csr_2511 = _RAND_2511[31:0];
  _RAND_2512 = {1{`RANDOM}};
  reg_csr_2512 = _RAND_2512[31:0];
  _RAND_2513 = {1{`RANDOM}};
  reg_csr_2513 = _RAND_2513[31:0];
  _RAND_2514 = {1{`RANDOM}};
  reg_csr_2514 = _RAND_2514[31:0];
  _RAND_2515 = {1{`RANDOM}};
  reg_csr_2515 = _RAND_2515[31:0];
  _RAND_2516 = {1{`RANDOM}};
  reg_csr_2516 = _RAND_2516[31:0];
  _RAND_2517 = {1{`RANDOM}};
  reg_csr_2517 = _RAND_2517[31:0];
  _RAND_2518 = {1{`RANDOM}};
  reg_csr_2518 = _RAND_2518[31:0];
  _RAND_2519 = {1{`RANDOM}};
  reg_csr_2519 = _RAND_2519[31:0];
  _RAND_2520 = {1{`RANDOM}};
  reg_csr_2520 = _RAND_2520[31:0];
  _RAND_2521 = {1{`RANDOM}};
  reg_csr_2521 = _RAND_2521[31:0];
  _RAND_2522 = {1{`RANDOM}};
  reg_csr_2522 = _RAND_2522[31:0];
  _RAND_2523 = {1{`RANDOM}};
  reg_csr_2523 = _RAND_2523[31:0];
  _RAND_2524 = {1{`RANDOM}};
  reg_csr_2524 = _RAND_2524[31:0];
  _RAND_2525 = {1{`RANDOM}};
  reg_csr_2525 = _RAND_2525[31:0];
  _RAND_2526 = {1{`RANDOM}};
  reg_csr_2526 = _RAND_2526[31:0];
  _RAND_2527 = {1{`RANDOM}};
  reg_csr_2527 = _RAND_2527[31:0];
  _RAND_2528 = {1{`RANDOM}};
  reg_csr_2528 = _RAND_2528[31:0];
  _RAND_2529 = {1{`RANDOM}};
  reg_csr_2529 = _RAND_2529[31:0];
  _RAND_2530 = {1{`RANDOM}};
  reg_csr_2530 = _RAND_2530[31:0];
  _RAND_2531 = {1{`RANDOM}};
  reg_csr_2531 = _RAND_2531[31:0];
  _RAND_2532 = {1{`RANDOM}};
  reg_csr_2532 = _RAND_2532[31:0];
  _RAND_2533 = {1{`RANDOM}};
  reg_csr_2533 = _RAND_2533[31:0];
  _RAND_2534 = {1{`RANDOM}};
  reg_csr_2534 = _RAND_2534[31:0];
  _RAND_2535 = {1{`RANDOM}};
  reg_csr_2535 = _RAND_2535[31:0];
  _RAND_2536 = {1{`RANDOM}};
  reg_csr_2536 = _RAND_2536[31:0];
  _RAND_2537 = {1{`RANDOM}};
  reg_csr_2537 = _RAND_2537[31:0];
  _RAND_2538 = {1{`RANDOM}};
  reg_csr_2538 = _RAND_2538[31:0];
  _RAND_2539 = {1{`RANDOM}};
  reg_csr_2539 = _RAND_2539[31:0];
  _RAND_2540 = {1{`RANDOM}};
  reg_csr_2540 = _RAND_2540[31:0];
  _RAND_2541 = {1{`RANDOM}};
  reg_csr_2541 = _RAND_2541[31:0];
  _RAND_2542 = {1{`RANDOM}};
  reg_csr_2542 = _RAND_2542[31:0];
  _RAND_2543 = {1{`RANDOM}};
  reg_csr_2543 = _RAND_2543[31:0];
  _RAND_2544 = {1{`RANDOM}};
  reg_csr_2544 = _RAND_2544[31:0];
  _RAND_2545 = {1{`RANDOM}};
  reg_csr_2545 = _RAND_2545[31:0];
  _RAND_2546 = {1{`RANDOM}};
  reg_csr_2546 = _RAND_2546[31:0];
  _RAND_2547 = {1{`RANDOM}};
  reg_csr_2547 = _RAND_2547[31:0];
  _RAND_2548 = {1{`RANDOM}};
  reg_csr_2548 = _RAND_2548[31:0];
  _RAND_2549 = {1{`RANDOM}};
  reg_csr_2549 = _RAND_2549[31:0];
  _RAND_2550 = {1{`RANDOM}};
  reg_csr_2550 = _RAND_2550[31:0];
  _RAND_2551 = {1{`RANDOM}};
  reg_csr_2551 = _RAND_2551[31:0];
  _RAND_2552 = {1{`RANDOM}};
  reg_csr_2552 = _RAND_2552[31:0];
  _RAND_2553 = {1{`RANDOM}};
  reg_csr_2553 = _RAND_2553[31:0];
  _RAND_2554 = {1{`RANDOM}};
  reg_csr_2554 = _RAND_2554[31:0];
  _RAND_2555 = {1{`RANDOM}};
  reg_csr_2555 = _RAND_2555[31:0];
  _RAND_2556 = {1{`RANDOM}};
  reg_csr_2556 = _RAND_2556[31:0];
  _RAND_2557 = {1{`RANDOM}};
  reg_csr_2557 = _RAND_2557[31:0];
  _RAND_2558 = {1{`RANDOM}};
  reg_csr_2558 = _RAND_2558[31:0];
  _RAND_2559 = {1{`RANDOM}};
  reg_csr_2559 = _RAND_2559[31:0];
  _RAND_2560 = {1{`RANDOM}};
  reg_csr_2560 = _RAND_2560[31:0];
  _RAND_2561 = {1{`RANDOM}};
  reg_csr_2561 = _RAND_2561[31:0];
  _RAND_2562 = {1{`RANDOM}};
  reg_csr_2562 = _RAND_2562[31:0];
  _RAND_2563 = {1{`RANDOM}};
  reg_csr_2563 = _RAND_2563[31:0];
  _RAND_2564 = {1{`RANDOM}};
  reg_csr_2564 = _RAND_2564[31:0];
  _RAND_2565 = {1{`RANDOM}};
  reg_csr_2565 = _RAND_2565[31:0];
  _RAND_2566 = {1{`RANDOM}};
  reg_csr_2566 = _RAND_2566[31:0];
  _RAND_2567 = {1{`RANDOM}};
  reg_csr_2567 = _RAND_2567[31:0];
  _RAND_2568 = {1{`RANDOM}};
  reg_csr_2568 = _RAND_2568[31:0];
  _RAND_2569 = {1{`RANDOM}};
  reg_csr_2569 = _RAND_2569[31:0];
  _RAND_2570 = {1{`RANDOM}};
  reg_csr_2570 = _RAND_2570[31:0];
  _RAND_2571 = {1{`RANDOM}};
  reg_csr_2571 = _RAND_2571[31:0];
  _RAND_2572 = {1{`RANDOM}};
  reg_csr_2572 = _RAND_2572[31:0];
  _RAND_2573 = {1{`RANDOM}};
  reg_csr_2573 = _RAND_2573[31:0];
  _RAND_2574 = {1{`RANDOM}};
  reg_csr_2574 = _RAND_2574[31:0];
  _RAND_2575 = {1{`RANDOM}};
  reg_csr_2575 = _RAND_2575[31:0];
  _RAND_2576 = {1{`RANDOM}};
  reg_csr_2576 = _RAND_2576[31:0];
  _RAND_2577 = {1{`RANDOM}};
  reg_csr_2577 = _RAND_2577[31:0];
  _RAND_2578 = {1{`RANDOM}};
  reg_csr_2578 = _RAND_2578[31:0];
  _RAND_2579 = {1{`RANDOM}};
  reg_csr_2579 = _RAND_2579[31:0];
  _RAND_2580 = {1{`RANDOM}};
  reg_csr_2580 = _RAND_2580[31:0];
  _RAND_2581 = {1{`RANDOM}};
  reg_csr_2581 = _RAND_2581[31:0];
  _RAND_2582 = {1{`RANDOM}};
  reg_csr_2582 = _RAND_2582[31:0];
  _RAND_2583 = {1{`RANDOM}};
  reg_csr_2583 = _RAND_2583[31:0];
  _RAND_2584 = {1{`RANDOM}};
  reg_csr_2584 = _RAND_2584[31:0];
  _RAND_2585 = {1{`RANDOM}};
  reg_csr_2585 = _RAND_2585[31:0];
  _RAND_2586 = {1{`RANDOM}};
  reg_csr_2586 = _RAND_2586[31:0];
  _RAND_2587 = {1{`RANDOM}};
  reg_csr_2587 = _RAND_2587[31:0];
  _RAND_2588 = {1{`RANDOM}};
  reg_csr_2588 = _RAND_2588[31:0];
  _RAND_2589 = {1{`RANDOM}};
  reg_csr_2589 = _RAND_2589[31:0];
  _RAND_2590 = {1{`RANDOM}};
  reg_csr_2590 = _RAND_2590[31:0];
  _RAND_2591 = {1{`RANDOM}};
  reg_csr_2591 = _RAND_2591[31:0];
  _RAND_2592 = {1{`RANDOM}};
  reg_csr_2592 = _RAND_2592[31:0];
  _RAND_2593 = {1{`RANDOM}};
  reg_csr_2593 = _RAND_2593[31:0];
  _RAND_2594 = {1{`RANDOM}};
  reg_csr_2594 = _RAND_2594[31:0];
  _RAND_2595 = {1{`RANDOM}};
  reg_csr_2595 = _RAND_2595[31:0];
  _RAND_2596 = {1{`RANDOM}};
  reg_csr_2596 = _RAND_2596[31:0];
  _RAND_2597 = {1{`RANDOM}};
  reg_csr_2597 = _RAND_2597[31:0];
  _RAND_2598 = {1{`RANDOM}};
  reg_csr_2598 = _RAND_2598[31:0];
  _RAND_2599 = {1{`RANDOM}};
  reg_csr_2599 = _RAND_2599[31:0];
  _RAND_2600 = {1{`RANDOM}};
  reg_csr_2600 = _RAND_2600[31:0];
  _RAND_2601 = {1{`RANDOM}};
  reg_csr_2601 = _RAND_2601[31:0];
  _RAND_2602 = {1{`RANDOM}};
  reg_csr_2602 = _RAND_2602[31:0];
  _RAND_2603 = {1{`RANDOM}};
  reg_csr_2603 = _RAND_2603[31:0];
  _RAND_2604 = {1{`RANDOM}};
  reg_csr_2604 = _RAND_2604[31:0];
  _RAND_2605 = {1{`RANDOM}};
  reg_csr_2605 = _RAND_2605[31:0];
  _RAND_2606 = {1{`RANDOM}};
  reg_csr_2606 = _RAND_2606[31:0];
  _RAND_2607 = {1{`RANDOM}};
  reg_csr_2607 = _RAND_2607[31:0];
  _RAND_2608 = {1{`RANDOM}};
  reg_csr_2608 = _RAND_2608[31:0];
  _RAND_2609 = {1{`RANDOM}};
  reg_csr_2609 = _RAND_2609[31:0];
  _RAND_2610 = {1{`RANDOM}};
  reg_csr_2610 = _RAND_2610[31:0];
  _RAND_2611 = {1{`RANDOM}};
  reg_csr_2611 = _RAND_2611[31:0];
  _RAND_2612 = {1{`RANDOM}};
  reg_csr_2612 = _RAND_2612[31:0];
  _RAND_2613 = {1{`RANDOM}};
  reg_csr_2613 = _RAND_2613[31:0];
  _RAND_2614 = {1{`RANDOM}};
  reg_csr_2614 = _RAND_2614[31:0];
  _RAND_2615 = {1{`RANDOM}};
  reg_csr_2615 = _RAND_2615[31:0];
  _RAND_2616 = {1{`RANDOM}};
  reg_csr_2616 = _RAND_2616[31:0];
  _RAND_2617 = {1{`RANDOM}};
  reg_csr_2617 = _RAND_2617[31:0];
  _RAND_2618 = {1{`RANDOM}};
  reg_csr_2618 = _RAND_2618[31:0];
  _RAND_2619 = {1{`RANDOM}};
  reg_csr_2619 = _RAND_2619[31:0];
  _RAND_2620 = {1{`RANDOM}};
  reg_csr_2620 = _RAND_2620[31:0];
  _RAND_2621 = {1{`RANDOM}};
  reg_csr_2621 = _RAND_2621[31:0];
  _RAND_2622 = {1{`RANDOM}};
  reg_csr_2622 = _RAND_2622[31:0];
  _RAND_2623 = {1{`RANDOM}};
  reg_csr_2623 = _RAND_2623[31:0];
  _RAND_2624 = {1{`RANDOM}};
  reg_csr_2624 = _RAND_2624[31:0];
  _RAND_2625 = {1{`RANDOM}};
  reg_csr_2625 = _RAND_2625[31:0];
  _RAND_2626 = {1{`RANDOM}};
  reg_csr_2626 = _RAND_2626[31:0];
  _RAND_2627 = {1{`RANDOM}};
  reg_csr_2627 = _RAND_2627[31:0];
  _RAND_2628 = {1{`RANDOM}};
  reg_csr_2628 = _RAND_2628[31:0];
  _RAND_2629 = {1{`RANDOM}};
  reg_csr_2629 = _RAND_2629[31:0];
  _RAND_2630 = {1{`RANDOM}};
  reg_csr_2630 = _RAND_2630[31:0];
  _RAND_2631 = {1{`RANDOM}};
  reg_csr_2631 = _RAND_2631[31:0];
  _RAND_2632 = {1{`RANDOM}};
  reg_csr_2632 = _RAND_2632[31:0];
  _RAND_2633 = {1{`RANDOM}};
  reg_csr_2633 = _RAND_2633[31:0];
  _RAND_2634 = {1{`RANDOM}};
  reg_csr_2634 = _RAND_2634[31:0];
  _RAND_2635 = {1{`RANDOM}};
  reg_csr_2635 = _RAND_2635[31:0];
  _RAND_2636 = {1{`RANDOM}};
  reg_csr_2636 = _RAND_2636[31:0];
  _RAND_2637 = {1{`RANDOM}};
  reg_csr_2637 = _RAND_2637[31:0];
  _RAND_2638 = {1{`RANDOM}};
  reg_csr_2638 = _RAND_2638[31:0];
  _RAND_2639 = {1{`RANDOM}};
  reg_csr_2639 = _RAND_2639[31:0];
  _RAND_2640 = {1{`RANDOM}};
  reg_csr_2640 = _RAND_2640[31:0];
  _RAND_2641 = {1{`RANDOM}};
  reg_csr_2641 = _RAND_2641[31:0];
  _RAND_2642 = {1{`RANDOM}};
  reg_csr_2642 = _RAND_2642[31:0];
  _RAND_2643 = {1{`RANDOM}};
  reg_csr_2643 = _RAND_2643[31:0];
  _RAND_2644 = {1{`RANDOM}};
  reg_csr_2644 = _RAND_2644[31:0];
  _RAND_2645 = {1{`RANDOM}};
  reg_csr_2645 = _RAND_2645[31:0];
  _RAND_2646 = {1{`RANDOM}};
  reg_csr_2646 = _RAND_2646[31:0];
  _RAND_2647 = {1{`RANDOM}};
  reg_csr_2647 = _RAND_2647[31:0];
  _RAND_2648 = {1{`RANDOM}};
  reg_csr_2648 = _RAND_2648[31:0];
  _RAND_2649 = {1{`RANDOM}};
  reg_csr_2649 = _RAND_2649[31:0];
  _RAND_2650 = {1{`RANDOM}};
  reg_csr_2650 = _RAND_2650[31:0];
  _RAND_2651 = {1{`RANDOM}};
  reg_csr_2651 = _RAND_2651[31:0];
  _RAND_2652 = {1{`RANDOM}};
  reg_csr_2652 = _RAND_2652[31:0];
  _RAND_2653 = {1{`RANDOM}};
  reg_csr_2653 = _RAND_2653[31:0];
  _RAND_2654 = {1{`RANDOM}};
  reg_csr_2654 = _RAND_2654[31:0];
  _RAND_2655 = {1{`RANDOM}};
  reg_csr_2655 = _RAND_2655[31:0];
  _RAND_2656 = {1{`RANDOM}};
  reg_csr_2656 = _RAND_2656[31:0];
  _RAND_2657 = {1{`RANDOM}};
  reg_csr_2657 = _RAND_2657[31:0];
  _RAND_2658 = {1{`RANDOM}};
  reg_csr_2658 = _RAND_2658[31:0];
  _RAND_2659 = {1{`RANDOM}};
  reg_csr_2659 = _RAND_2659[31:0];
  _RAND_2660 = {1{`RANDOM}};
  reg_csr_2660 = _RAND_2660[31:0];
  _RAND_2661 = {1{`RANDOM}};
  reg_csr_2661 = _RAND_2661[31:0];
  _RAND_2662 = {1{`RANDOM}};
  reg_csr_2662 = _RAND_2662[31:0];
  _RAND_2663 = {1{`RANDOM}};
  reg_csr_2663 = _RAND_2663[31:0];
  _RAND_2664 = {1{`RANDOM}};
  reg_csr_2664 = _RAND_2664[31:0];
  _RAND_2665 = {1{`RANDOM}};
  reg_csr_2665 = _RAND_2665[31:0];
  _RAND_2666 = {1{`RANDOM}};
  reg_csr_2666 = _RAND_2666[31:0];
  _RAND_2667 = {1{`RANDOM}};
  reg_csr_2667 = _RAND_2667[31:0];
  _RAND_2668 = {1{`RANDOM}};
  reg_csr_2668 = _RAND_2668[31:0];
  _RAND_2669 = {1{`RANDOM}};
  reg_csr_2669 = _RAND_2669[31:0];
  _RAND_2670 = {1{`RANDOM}};
  reg_csr_2670 = _RAND_2670[31:0];
  _RAND_2671 = {1{`RANDOM}};
  reg_csr_2671 = _RAND_2671[31:0];
  _RAND_2672 = {1{`RANDOM}};
  reg_csr_2672 = _RAND_2672[31:0];
  _RAND_2673 = {1{`RANDOM}};
  reg_csr_2673 = _RAND_2673[31:0];
  _RAND_2674 = {1{`RANDOM}};
  reg_csr_2674 = _RAND_2674[31:0];
  _RAND_2675 = {1{`RANDOM}};
  reg_csr_2675 = _RAND_2675[31:0];
  _RAND_2676 = {1{`RANDOM}};
  reg_csr_2676 = _RAND_2676[31:0];
  _RAND_2677 = {1{`RANDOM}};
  reg_csr_2677 = _RAND_2677[31:0];
  _RAND_2678 = {1{`RANDOM}};
  reg_csr_2678 = _RAND_2678[31:0];
  _RAND_2679 = {1{`RANDOM}};
  reg_csr_2679 = _RAND_2679[31:0];
  _RAND_2680 = {1{`RANDOM}};
  reg_csr_2680 = _RAND_2680[31:0];
  _RAND_2681 = {1{`RANDOM}};
  reg_csr_2681 = _RAND_2681[31:0];
  _RAND_2682 = {1{`RANDOM}};
  reg_csr_2682 = _RAND_2682[31:0];
  _RAND_2683 = {1{`RANDOM}};
  reg_csr_2683 = _RAND_2683[31:0];
  _RAND_2684 = {1{`RANDOM}};
  reg_csr_2684 = _RAND_2684[31:0];
  _RAND_2685 = {1{`RANDOM}};
  reg_csr_2685 = _RAND_2685[31:0];
  _RAND_2686 = {1{`RANDOM}};
  reg_csr_2686 = _RAND_2686[31:0];
  _RAND_2687 = {1{`RANDOM}};
  reg_csr_2687 = _RAND_2687[31:0];
  _RAND_2688 = {1{`RANDOM}};
  reg_csr_2688 = _RAND_2688[31:0];
  _RAND_2689 = {1{`RANDOM}};
  reg_csr_2689 = _RAND_2689[31:0];
  _RAND_2690 = {1{`RANDOM}};
  reg_csr_2690 = _RAND_2690[31:0];
  _RAND_2691 = {1{`RANDOM}};
  reg_csr_2691 = _RAND_2691[31:0];
  _RAND_2692 = {1{`RANDOM}};
  reg_csr_2692 = _RAND_2692[31:0];
  _RAND_2693 = {1{`RANDOM}};
  reg_csr_2693 = _RAND_2693[31:0];
  _RAND_2694 = {1{`RANDOM}};
  reg_csr_2694 = _RAND_2694[31:0];
  _RAND_2695 = {1{`RANDOM}};
  reg_csr_2695 = _RAND_2695[31:0];
  _RAND_2696 = {1{`RANDOM}};
  reg_csr_2696 = _RAND_2696[31:0];
  _RAND_2697 = {1{`RANDOM}};
  reg_csr_2697 = _RAND_2697[31:0];
  _RAND_2698 = {1{`RANDOM}};
  reg_csr_2698 = _RAND_2698[31:0];
  _RAND_2699 = {1{`RANDOM}};
  reg_csr_2699 = _RAND_2699[31:0];
  _RAND_2700 = {1{`RANDOM}};
  reg_csr_2700 = _RAND_2700[31:0];
  _RAND_2701 = {1{`RANDOM}};
  reg_csr_2701 = _RAND_2701[31:0];
  _RAND_2702 = {1{`RANDOM}};
  reg_csr_2702 = _RAND_2702[31:0];
  _RAND_2703 = {1{`RANDOM}};
  reg_csr_2703 = _RAND_2703[31:0];
  _RAND_2704 = {1{`RANDOM}};
  reg_csr_2704 = _RAND_2704[31:0];
  _RAND_2705 = {1{`RANDOM}};
  reg_csr_2705 = _RAND_2705[31:0];
  _RAND_2706 = {1{`RANDOM}};
  reg_csr_2706 = _RAND_2706[31:0];
  _RAND_2707 = {1{`RANDOM}};
  reg_csr_2707 = _RAND_2707[31:0];
  _RAND_2708 = {1{`RANDOM}};
  reg_csr_2708 = _RAND_2708[31:0];
  _RAND_2709 = {1{`RANDOM}};
  reg_csr_2709 = _RAND_2709[31:0];
  _RAND_2710 = {1{`RANDOM}};
  reg_csr_2710 = _RAND_2710[31:0];
  _RAND_2711 = {1{`RANDOM}};
  reg_csr_2711 = _RAND_2711[31:0];
  _RAND_2712 = {1{`RANDOM}};
  reg_csr_2712 = _RAND_2712[31:0];
  _RAND_2713 = {1{`RANDOM}};
  reg_csr_2713 = _RAND_2713[31:0];
  _RAND_2714 = {1{`RANDOM}};
  reg_csr_2714 = _RAND_2714[31:0];
  _RAND_2715 = {1{`RANDOM}};
  reg_csr_2715 = _RAND_2715[31:0];
  _RAND_2716 = {1{`RANDOM}};
  reg_csr_2716 = _RAND_2716[31:0];
  _RAND_2717 = {1{`RANDOM}};
  reg_csr_2717 = _RAND_2717[31:0];
  _RAND_2718 = {1{`RANDOM}};
  reg_csr_2718 = _RAND_2718[31:0];
  _RAND_2719 = {1{`RANDOM}};
  reg_csr_2719 = _RAND_2719[31:0];
  _RAND_2720 = {1{`RANDOM}};
  reg_csr_2720 = _RAND_2720[31:0];
  _RAND_2721 = {1{`RANDOM}};
  reg_csr_2721 = _RAND_2721[31:0];
  _RAND_2722 = {1{`RANDOM}};
  reg_csr_2722 = _RAND_2722[31:0];
  _RAND_2723 = {1{`RANDOM}};
  reg_csr_2723 = _RAND_2723[31:0];
  _RAND_2724 = {1{`RANDOM}};
  reg_csr_2724 = _RAND_2724[31:0];
  _RAND_2725 = {1{`RANDOM}};
  reg_csr_2725 = _RAND_2725[31:0];
  _RAND_2726 = {1{`RANDOM}};
  reg_csr_2726 = _RAND_2726[31:0];
  _RAND_2727 = {1{`RANDOM}};
  reg_csr_2727 = _RAND_2727[31:0];
  _RAND_2728 = {1{`RANDOM}};
  reg_csr_2728 = _RAND_2728[31:0];
  _RAND_2729 = {1{`RANDOM}};
  reg_csr_2729 = _RAND_2729[31:0];
  _RAND_2730 = {1{`RANDOM}};
  reg_csr_2730 = _RAND_2730[31:0];
  _RAND_2731 = {1{`RANDOM}};
  reg_csr_2731 = _RAND_2731[31:0];
  _RAND_2732 = {1{`RANDOM}};
  reg_csr_2732 = _RAND_2732[31:0];
  _RAND_2733 = {1{`RANDOM}};
  reg_csr_2733 = _RAND_2733[31:0];
  _RAND_2734 = {1{`RANDOM}};
  reg_csr_2734 = _RAND_2734[31:0];
  _RAND_2735 = {1{`RANDOM}};
  reg_csr_2735 = _RAND_2735[31:0];
  _RAND_2736 = {1{`RANDOM}};
  reg_csr_2736 = _RAND_2736[31:0];
  _RAND_2737 = {1{`RANDOM}};
  reg_csr_2737 = _RAND_2737[31:0];
  _RAND_2738 = {1{`RANDOM}};
  reg_csr_2738 = _RAND_2738[31:0];
  _RAND_2739 = {1{`RANDOM}};
  reg_csr_2739 = _RAND_2739[31:0];
  _RAND_2740 = {1{`RANDOM}};
  reg_csr_2740 = _RAND_2740[31:0];
  _RAND_2741 = {1{`RANDOM}};
  reg_csr_2741 = _RAND_2741[31:0];
  _RAND_2742 = {1{`RANDOM}};
  reg_csr_2742 = _RAND_2742[31:0];
  _RAND_2743 = {1{`RANDOM}};
  reg_csr_2743 = _RAND_2743[31:0];
  _RAND_2744 = {1{`RANDOM}};
  reg_csr_2744 = _RAND_2744[31:0];
  _RAND_2745 = {1{`RANDOM}};
  reg_csr_2745 = _RAND_2745[31:0];
  _RAND_2746 = {1{`RANDOM}};
  reg_csr_2746 = _RAND_2746[31:0];
  _RAND_2747 = {1{`RANDOM}};
  reg_csr_2747 = _RAND_2747[31:0];
  _RAND_2748 = {1{`RANDOM}};
  reg_csr_2748 = _RAND_2748[31:0];
  _RAND_2749 = {1{`RANDOM}};
  reg_csr_2749 = _RAND_2749[31:0];
  _RAND_2750 = {1{`RANDOM}};
  reg_csr_2750 = _RAND_2750[31:0];
  _RAND_2751 = {1{`RANDOM}};
  reg_csr_2751 = _RAND_2751[31:0];
  _RAND_2752 = {1{`RANDOM}};
  reg_csr_2752 = _RAND_2752[31:0];
  _RAND_2753 = {1{`RANDOM}};
  reg_csr_2753 = _RAND_2753[31:0];
  _RAND_2754 = {1{`RANDOM}};
  reg_csr_2754 = _RAND_2754[31:0];
  _RAND_2755 = {1{`RANDOM}};
  reg_csr_2755 = _RAND_2755[31:0];
  _RAND_2756 = {1{`RANDOM}};
  reg_csr_2756 = _RAND_2756[31:0];
  _RAND_2757 = {1{`RANDOM}};
  reg_csr_2757 = _RAND_2757[31:0];
  _RAND_2758 = {1{`RANDOM}};
  reg_csr_2758 = _RAND_2758[31:0];
  _RAND_2759 = {1{`RANDOM}};
  reg_csr_2759 = _RAND_2759[31:0];
  _RAND_2760 = {1{`RANDOM}};
  reg_csr_2760 = _RAND_2760[31:0];
  _RAND_2761 = {1{`RANDOM}};
  reg_csr_2761 = _RAND_2761[31:0];
  _RAND_2762 = {1{`RANDOM}};
  reg_csr_2762 = _RAND_2762[31:0];
  _RAND_2763 = {1{`RANDOM}};
  reg_csr_2763 = _RAND_2763[31:0];
  _RAND_2764 = {1{`RANDOM}};
  reg_csr_2764 = _RAND_2764[31:0];
  _RAND_2765 = {1{`RANDOM}};
  reg_csr_2765 = _RAND_2765[31:0];
  _RAND_2766 = {1{`RANDOM}};
  reg_csr_2766 = _RAND_2766[31:0];
  _RAND_2767 = {1{`RANDOM}};
  reg_csr_2767 = _RAND_2767[31:0];
  _RAND_2768 = {1{`RANDOM}};
  reg_csr_2768 = _RAND_2768[31:0];
  _RAND_2769 = {1{`RANDOM}};
  reg_csr_2769 = _RAND_2769[31:0];
  _RAND_2770 = {1{`RANDOM}};
  reg_csr_2770 = _RAND_2770[31:0];
  _RAND_2771 = {1{`RANDOM}};
  reg_csr_2771 = _RAND_2771[31:0];
  _RAND_2772 = {1{`RANDOM}};
  reg_csr_2772 = _RAND_2772[31:0];
  _RAND_2773 = {1{`RANDOM}};
  reg_csr_2773 = _RAND_2773[31:0];
  _RAND_2774 = {1{`RANDOM}};
  reg_csr_2774 = _RAND_2774[31:0];
  _RAND_2775 = {1{`RANDOM}};
  reg_csr_2775 = _RAND_2775[31:0];
  _RAND_2776 = {1{`RANDOM}};
  reg_csr_2776 = _RAND_2776[31:0];
  _RAND_2777 = {1{`RANDOM}};
  reg_csr_2777 = _RAND_2777[31:0];
  _RAND_2778 = {1{`RANDOM}};
  reg_csr_2778 = _RAND_2778[31:0];
  _RAND_2779 = {1{`RANDOM}};
  reg_csr_2779 = _RAND_2779[31:0];
  _RAND_2780 = {1{`RANDOM}};
  reg_csr_2780 = _RAND_2780[31:0];
  _RAND_2781 = {1{`RANDOM}};
  reg_csr_2781 = _RAND_2781[31:0];
  _RAND_2782 = {1{`RANDOM}};
  reg_csr_2782 = _RAND_2782[31:0];
  _RAND_2783 = {1{`RANDOM}};
  reg_csr_2783 = _RAND_2783[31:0];
  _RAND_2784 = {1{`RANDOM}};
  reg_csr_2784 = _RAND_2784[31:0];
  _RAND_2785 = {1{`RANDOM}};
  reg_csr_2785 = _RAND_2785[31:0];
  _RAND_2786 = {1{`RANDOM}};
  reg_csr_2786 = _RAND_2786[31:0];
  _RAND_2787 = {1{`RANDOM}};
  reg_csr_2787 = _RAND_2787[31:0];
  _RAND_2788 = {1{`RANDOM}};
  reg_csr_2788 = _RAND_2788[31:0];
  _RAND_2789 = {1{`RANDOM}};
  reg_csr_2789 = _RAND_2789[31:0];
  _RAND_2790 = {1{`RANDOM}};
  reg_csr_2790 = _RAND_2790[31:0];
  _RAND_2791 = {1{`RANDOM}};
  reg_csr_2791 = _RAND_2791[31:0];
  _RAND_2792 = {1{`RANDOM}};
  reg_csr_2792 = _RAND_2792[31:0];
  _RAND_2793 = {1{`RANDOM}};
  reg_csr_2793 = _RAND_2793[31:0];
  _RAND_2794 = {1{`RANDOM}};
  reg_csr_2794 = _RAND_2794[31:0];
  _RAND_2795 = {1{`RANDOM}};
  reg_csr_2795 = _RAND_2795[31:0];
  _RAND_2796 = {1{`RANDOM}};
  reg_csr_2796 = _RAND_2796[31:0];
  _RAND_2797 = {1{`RANDOM}};
  reg_csr_2797 = _RAND_2797[31:0];
  _RAND_2798 = {1{`RANDOM}};
  reg_csr_2798 = _RAND_2798[31:0];
  _RAND_2799 = {1{`RANDOM}};
  reg_csr_2799 = _RAND_2799[31:0];
  _RAND_2800 = {1{`RANDOM}};
  reg_csr_2800 = _RAND_2800[31:0];
  _RAND_2801 = {1{`RANDOM}};
  reg_csr_2801 = _RAND_2801[31:0];
  _RAND_2802 = {1{`RANDOM}};
  reg_csr_2802 = _RAND_2802[31:0];
  _RAND_2803 = {1{`RANDOM}};
  reg_csr_2803 = _RAND_2803[31:0];
  _RAND_2804 = {1{`RANDOM}};
  reg_csr_2804 = _RAND_2804[31:0];
  _RAND_2805 = {1{`RANDOM}};
  reg_csr_2805 = _RAND_2805[31:0];
  _RAND_2806 = {1{`RANDOM}};
  reg_csr_2806 = _RAND_2806[31:0];
  _RAND_2807 = {1{`RANDOM}};
  reg_csr_2807 = _RAND_2807[31:0];
  _RAND_2808 = {1{`RANDOM}};
  reg_csr_2808 = _RAND_2808[31:0];
  _RAND_2809 = {1{`RANDOM}};
  reg_csr_2809 = _RAND_2809[31:0];
  _RAND_2810 = {1{`RANDOM}};
  reg_csr_2810 = _RAND_2810[31:0];
  _RAND_2811 = {1{`RANDOM}};
  reg_csr_2811 = _RAND_2811[31:0];
  _RAND_2812 = {1{`RANDOM}};
  reg_csr_2812 = _RAND_2812[31:0];
  _RAND_2813 = {1{`RANDOM}};
  reg_csr_2813 = _RAND_2813[31:0];
  _RAND_2814 = {1{`RANDOM}};
  reg_csr_2814 = _RAND_2814[31:0];
  _RAND_2815 = {1{`RANDOM}};
  reg_csr_2815 = _RAND_2815[31:0];
  _RAND_2816 = {1{`RANDOM}};
  reg_csr_2816 = _RAND_2816[31:0];
  _RAND_2817 = {1{`RANDOM}};
  reg_csr_2817 = _RAND_2817[31:0];
  _RAND_2818 = {1{`RANDOM}};
  reg_csr_2818 = _RAND_2818[31:0];
  _RAND_2819 = {1{`RANDOM}};
  reg_csr_2819 = _RAND_2819[31:0];
  _RAND_2820 = {1{`RANDOM}};
  reg_csr_2820 = _RAND_2820[31:0];
  _RAND_2821 = {1{`RANDOM}};
  reg_csr_2821 = _RAND_2821[31:0];
  _RAND_2822 = {1{`RANDOM}};
  reg_csr_2822 = _RAND_2822[31:0];
  _RAND_2823 = {1{`RANDOM}};
  reg_csr_2823 = _RAND_2823[31:0];
  _RAND_2824 = {1{`RANDOM}};
  reg_csr_2824 = _RAND_2824[31:0];
  _RAND_2825 = {1{`RANDOM}};
  reg_csr_2825 = _RAND_2825[31:0];
  _RAND_2826 = {1{`RANDOM}};
  reg_csr_2826 = _RAND_2826[31:0];
  _RAND_2827 = {1{`RANDOM}};
  reg_csr_2827 = _RAND_2827[31:0];
  _RAND_2828 = {1{`RANDOM}};
  reg_csr_2828 = _RAND_2828[31:0];
  _RAND_2829 = {1{`RANDOM}};
  reg_csr_2829 = _RAND_2829[31:0];
  _RAND_2830 = {1{`RANDOM}};
  reg_csr_2830 = _RAND_2830[31:0];
  _RAND_2831 = {1{`RANDOM}};
  reg_csr_2831 = _RAND_2831[31:0];
  _RAND_2832 = {1{`RANDOM}};
  reg_csr_2832 = _RAND_2832[31:0];
  _RAND_2833 = {1{`RANDOM}};
  reg_csr_2833 = _RAND_2833[31:0];
  _RAND_2834 = {1{`RANDOM}};
  reg_csr_2834 = _RAND_2834[31:0];
  _RAND_2835 = {1{`RANDOM}};
  reg_csr_2835 = _RAND_2835[31:0];
  _RAND_2836 = {1{`RANDOM}};
  reg_csr_2836 = _RAND_2836[31:0];
  _RAND_2837 = {1{`RANDOM}};
  reg_csr_2837 = _RAND_2837[31:0];
  _RAND_2838 = {1{`RANDOM}};
  reg_csr_2838 = _RAND_2838[31:0];
  _RAND_2839 = {1{`RANDOM}};
  reg_csr_2839 = _RAND_2839[31:0];
  _RAND_2840 = {1{`RANDOM}};
  reg_csr_2840 = _RAND_2840[31:0];
  _RAND_2841 = {1{`RANDOM}};
  reg_csr_2841 = _RAND_2841[31:0];
  _RAND_2842 = {1{`RANDOM}};
  reg_csr_2842 = _RAND_2842[31:0];
  _RAND_2843 = {1{`RANDOM}};
  reg_csr_2843 = _RAND_2843[31:0];
  _RAND_2844 = {1{`RANDOM}};
  reg_csr_2844 = _RAND_2844[31:0];
  _RAND_2845 = {1{`RANDOM}};
  reg_csr_2845 = _RAND_2845[31:0];
  _RAND_2846 = {1{`RANDOM}};
  reg_csr_2846 = _RAND_2846[31:0];
  _RAND_2847 = {1{`RANDOM}};
  reg_csr_2847 = _RAND_2847[31:0];
  _RAND_2848 = {1{`RANDOM}};
  reg_csr_2848 = _RAND_2848[31:0];
  _RAND_2849 = {1{`RANDOM}};
  reg_csr_2849 = _RAND_2849[31:0];
  _RAND_2850 = {1{`RANDOM}};
  reg_csr_2850 = _RAND_2850[31:0];
  _RAND_2851 = {1{`RANDOM}};
  reg_csr_2851 = _RAND_2851[31:0];
  _RAND_2852 = {1{`RANDOM}};
  reg_csr_2852 = _RAND_2852[31:0];
  _RAND_2853 = {1{`RANDOM}};
  reg_csr_2853 = _RAND_2853[31:0];
  _RAND_2854 = {1{`RANDOM}};
  reg_csr_2854 = _RAND_2854[31:0];
  _RAND_2855 = {1{`RANDOM}};
  reg_csr_2855 = _RAND_2855[31:0];
  _RAND_2856 = {1{`RANDOM}};
  reg_csr_2856 = _RAND_2856[31:0];
  _RAND_2857 = {1{`RANDOM}};
  reg_csr_2857 = _RAND_2857[31:0];
  _RAND_2858 = {1{`RANDOM}};
  reg_csr_2858 = _RAND_2858[31:0];
  _RAND_2859 = {1{`RANDOM}};
  reg_csr_2859 = _RAND_2859[31:0];
  _RAND_2860 = {1{`RANDOM}};
  reg_csr_2860 = _RAND_2860[31:0];
  _RAND_2861 = {1{`RANDOM}};
  reg_csr_2861 = _RAND_2861[31:0];
  _RAND_2862 = {1{`RANDOM}};
  reg_csr_2862 = _RAND_2862[31:0];
  _RAND_2863 = {1{`RANDOM}};
  reg_csr_2863 = _RAND_2863[31:0];
  _RAND_2864 = {1{`RANDOM}};
  reg_csr_2864 = _RAND_2864[31:0];
  _RAND_2865 = {1{`RANDOM}};
  reg_csr_2865 = _RAND_2865[31:0];
  _RAND_2866 = {1{`RANDOM}};
  reg_csr_2866 = _RAND_2866[31:0];
  _RAND_2867 = {1{`RANDOM}};
  reg_csr_2867 = _RAND_2867[31:0];
  _RAND_2868 = {1{`RANDOM}};
  reg_csr_2868 = _RAND_2868[31:0];
  _RAND_2869 = {1{`RANDOM}};
  reg_csr_2869 = _RAND_2869[31:0];
  _RAND_2870 = {1{`RANDOM}};
  reg_csr_2870 = _RAND_2870[31:0];
  _RAND_2871 = {1{`RANDOM}};
  reg_csr_2871 = _RAND_2871[31:0];
  _RAND_2872 = {1{`RANDOM}};
  reg_csr_2872 = _RAND_2872[31:0];
  _RAND_2873 = {1{`RANDOM}};
  reg_csr_2873 = _RAND_2873[31:0];
  _RAND_2874 = {1{`RANDOM}};
  reg_csr_2874 = _RAND_2874[31:0];
  _RAND_2875 = {1{`RANDOM}};
  reg_csr_2875 = _RAND_2875[31:0];
  _RAND_2876 = {1{`RANDOM}};
  reg_csr_2876 = _RAND_2876[31:0];
  _RAND_2877 = {1{`RANDOM}};
  reg_csr_2877 = _RAND_2877[31:0];
  _RAND_2878 = {1{`RANDOM}};
  reg_csr_2878 = _RAND_2878[31:0];
  _RAND_2879 = {1{`RANDOM}};
  reg_csr_2879 = _RAND_2879[31:0];
  _RAND_2880 = {1{`RANDOM}};
  reg_csr_2880 = _RAND_2880[31:0];
  _RAND_2881 = {1{`RANDOM}};
  reg_csr_2881 = _RAND_2881[31:0];
  _RAND_2882 = {1{`RANDOM}};
  reg_csr_2882 = _RAND_2882[31:0];
  _RAND_2883 = {1{`RANDOM}};
  reg_csr_2883 = _RAND_2883[31:0];
  _RAND_2884 = {1{`RANDOM}};
  reg_csr_2884 = _RAND_2884[31:0];
  _RAND_2885 = {1{`RANDOM}};
  reg_csr_2885 = _RAND_2885[31:0];
  _RAND_2886 = {1{`RANDOM}};
  reg_csr_2886 = _RAND_2886[31:0];
  _RAND_2887 = {1{`RANDOM}};
  reg_csr_2887 = _RAND_2887[31:0];
  _RAND_2888 = {1{`RANDOM}};
  reg_csr_2888 = _RAND_2888[31:0];
  _RAND_2889 = {1{`RANDOM}};
  reg_csr_2889 = _RAND_2889[31:0];
  _RAND_2890 = {1{`RANDOM}};
  reg_csr_2890 = _RAND_2890[31:0];
  _RAND_2891 = {1{`RANDOM}};
  reg_csr_2891 = _RAND_2891[31:0];
  _RAND_2892 = {1{`RANDOM}};
  reg_csr_2892 = _RAND_2892[31:0];
  _RAND_2893 = {1{`RANDOM}};
  reg_csr_2893 = _RAND_2893[31:0];
  _RAND_2894 = {1{`RANDOM}};
  reg_csr_2894 = _RAND_2894[31:0];
  _RAND_2895 = {1{`RANDOM}};
  reg_csr_2895 = _RAND_2895[31:0];
  _RAND_2896 = {1{`RANDOM}};
  reg_csr_2896 = _RAND_2896[31:0];
  _RAND_2897 = {1{`RANDOM}};
  reg_csr_2897 = _RAND_2897[31:0];
  _RAND_2898 = {1{`RANDOM}};
  reg_csr_2898 = _RAND_2898[31:0];
  _RAND_2899 = {1{`RANDOM}};
  reg_csr_2899 = _RAND_2899[31:0];
  _RAND_2900 = {1{`RANDOM}};
  reg_csr_2900 = _RAND_2900[31:0];
  _RAND_2901 = {1{`RANDOM}};
  reg_csr_2901 = _RAND_2901[31:0];
  _RAND_2902 = {1{`RANDOM}};
  reg_csr_2902 = _RAND_2902[31:0];
  _RAND_2903 = {1{`RANDOM}};
  reg_csr_2903 = _RAND_2903[31:0];
  _RAND_2904 = {1{`RANDOM}};
  reg_csr_2904 = _RAND_2904[31:0];
  _RAND_2905 = {1{`RANDOM}};
  reg_csr_2905 = _RAND_2905[31:0];
  _RAND_2906 = {1{`RANDOM}};
  reg_csr_2906 = _RAND_2906[31:0];
  _RAND_2907 = {1{`RANDOM}};
  reg_csr_2907 = _RAND_2907[31:0];
  _RAND_2908 = {1{`RANDOM}};
  reg_csr_2908 = _RAND_2908[31:0];
  _RAND_2909 = {1{`RANDOM}};
  reg_csr_2909 = _RAND_2909[31:0];
  _RAND_2910 = {1{`RANDOM}};
  reg_csr_2910 = _RAND_2910[31:0];
  _RAND_2911 = {1{`RANDOM}};
  reg_csr_2911 = _RAND_2911[31:0];
  _RAND_2912 = {1{`RANDOM}};
  reg_csr_2912 = _RAND_2912[31:0];
  _RAND_2913 = {1{`RANDOM}};
  reg_csr_2913 = _RAND_2913[31:0];
  _RAND_2914 = {1{`RANDOM}};
  reg_csr_2914 = _RAND_2914[31:0];
  _RAND_2915 = {1{`RANDOM}};
  reg_csr_2915 = _RAND_2915[31:0];
  _RAND_2916 = {1{`RANDOM}};
  reg_csr_2916 = _RAND_2916[31:0];
  _RAND_2917 = {1{`RANDOM}};
  reg_csr_2917 = _RAND_2917[31:0];
  _RAND_2918 = {1{`RANDOM}};
  reg_csr_2918 = _RAND_2918[31:0];
  _RAND_2919 = {1{`RANDOM}};
  reg_csr_2919 = _RAND_2919[31:0];
  _RAND_2920 = {1{`RANDOM}};
  reg_csr_2920 = _RAND_2920[31:0];
  _RAND_2921 = {1{`RANDOM}};
  reg_csr_2921 = _RAND_2921[31:0];
  _RAND_2922 = {1{`RANDOM}};
  reg_csr_2922 = _RAND_2922[31:0];
  _RAND_2923 = {1{`RANDOM}};
  reg_csr_2923 = _RAND_2923[31:0];
  _RAND_2924 = {1{`RANDOM}};
  reg_csr_2924 = _RAND_2924[31:0];
  _RAND_2925 = {1{`RANDOM}};
  reg_csr_2925 = _RAND_2925[31:0];
  _RAND_2926 = {1{`RANDOM}};
  reg_csr_2926 = _RAND_2926[31:0];
  _RAND_2927 = {1{`RANDOM}};
  reg_csr_2927 = _RAND_2927[31:0];
  _RAND_2928 = {1{`RANDOM}};
  reg_csr_2928 = _RAND_2928[31:0];
  _RAND_2929 = {1{`RANDOM}};
  reg_csr_2929 = _RAND_2929[31:0];
  _RAND_2930 = {1{`RANDOM}};
  reg_csr_2930 = _RAND_2930[31:0];
  _RAND_2931 = {1{`RANDOM}};
  reg_csr_2931 = _RAND_2931[31:0];
  _RAND_2932 = {1{`RANDOM}};
  reg_csr_2932 = _RAND_2932[31:0];
  _RAND_2933 = {1{`RANDOM}};
  reg_csr_2933 = _RAND_2933[31:0];
  _RAND_2934 = {1{`RANDOM}};
  reg_csr_2934 = _RAND_2934[31:0];
  _RAND_2935 = {1{`RANDOM}};
  reg_csr_2935 = _RAND_2935[31:0];
  _RAND_2936 = {1{`RANDOM}};
  reg_csr_2936 = _RAND_2936[31:0];
  _RAND_2937 = {1{`RANDOM}};
  reg_csr_2937 = _RAND_2937[31:0];
  _RAND_2938 = {1{`RANDOM}};
  reg_csr_2938 = _RAND_2938[31:0];
  _RAND_2939 = {1{`RANDOM}};
  reg_csr_2939 = _RAND_2939[31:0];
  _RAND_2940 = {1{`RANDOM}};
  reg_csr_2940 = _RAND_2940[31:0];
  _RAND_2941 = {1{`RANDOM}};
  reg_csr_2941 = _RAND_2941[31:0];
  _RAND_2942 = {1{`RANDOM}};
  reg_csr_2942 = _RAND_2942[31:0];
  _RAND_2943 = {1{`RANDOM}};
  reg_csr_2943 = _RAND_2943[31:0];
  _RAND_2944 = {1{`RANDOM}};
  reg_csr_2944 = _RAND_2944[31:0];
  _RAND_2945 = {1{`RANDOM}};
  reg_csr_2945 = _RAND_2945[31:0];
  _RAND_2946 = {1{`RANDOM}};
  reg_csr_2946 = _RAND_2946[31:0];
  _RAND_2947 = {1{`RANDOM}};
  reg_csr_2947 = _RAND_2947[31:0];
  _RAND_2948 = {1{`RANDOM}};
  reg_csr_2948 = _RAND_2948[31:0];
  _RAND_2949 = {1{`RANDOM}};
  reg_csr_2949 = _RAND_2949[31:0];
  _RAND_2950 = {1{`RANDOM}};
  reg_csr_2950 = _RAND_2950[31:0];
  _RAND_2951 = {1{`RANDOM}};
  reg_csr_2951 = _RAND_2951[31:0];
  _RAND_2952 = {1{`RANDOM}};
  reg_csr_2952 = _RAND_2952[31:0];
  _RAND_2953 = {1{`RANDOM}};
  reg_csr_2953 = _RAND_2953[31:0];
  _RAND_2954 = {1{`RANDOM}};
  reg_csr_2954 = _RAND_2954[31:0];
  _RAND_2955 = {1{`RANDOM}};
  reg_csr_2955 = _RAND_2955[31:0];
  _RAND_2956 = {1{`RANDOM}};
  reg_csr_2956 = _RAND_2956[31:0];
  _RAND_2957 = {1{`RANDOM}};
  reg_csr_2957 = _RAND_2957[31:0];
  _RAND_2958 = {1{`RANDOM}};
  reg_csr_2958 = _RAND_2958[31:0];
  _RAND_2959 = {1{`RANDOM}};
  reg_csr_2959 = _RAND_2959[31:0];
  _RAND_2960 = {1{`RANDOM}};
  reg_csr_2960 = _RAND_2960[31:0];
  _RAND_2961 = {1{`RANDOM}};
  reg_csr_2961 = _RAND_2961[31:0];
  _RAND_2962 = {1{`RANDOM}};
  reg_csr_2962 = _RAND_2962[31:0];
  _RAND_2963 = {1{`RANDOM}};
  reg_csr_2963 = _RAND_2963[31:0];
  _RAND_2964 = {1{`RANDOM}};
  reg_csr_2964 = _RAND_2964[31:0];
  _RAND_2965 = {1{`RANDOM}};
  reg_csr_2965 = _RAND_2965[31:0];
  _RAND_2966 = {1{`RANDOM}};
  reg_csr_2966 = _RAND_2966[31:0];
  _RAND_2967 = {1{`RANDOM}};
  reg_csr_2967 = _RAND_2967[31:0];
  _RAND_2968 = {1{`RANDOM}};
  reg_csr_2968 = _RAND_2968[31:0];
  _RAND_2969 = {1{`RANDOM}};
  reg_csr_2969 = _RAND_2969[31:0];
  _RAND_2970 = {1{`RANDOM}};
  reg_csr_2970 = _RAND_2970[31:0];
  _RAND_2971 = {1{`RANDOM}};
  reg_csr_2971 = _RAND_2971[31:0];
  _RAND_2972 = {1{`RANDOM}};
  reg_csr_2972 = _RAND_2972[31:0];
  _RAND_2973 = {1{`RANDOM}};
  reg_csr_2973 = _RAND_2973[31:0];
  _RAND_2974 = {1{`RANDOM}};
  reg_csr_2974 = _RAND_2974[31:0];
  _RAND_2975 = {1{`RANDOM}};
  reg_csr_2975 = _RAND_2975[31:0];
  _RAND_2976 = {1{`RANDOM}};
  reg_csr_2976 = _RAND_2976[31:0];
  _RAND_2977 = {1{`RANDOM}};
  reg_csr_2977 = _RAND_2977[31:0];
  _RAND_2978 = {1{`RANDOM}};
  reg_csr_2978 = _RAND_2978[31:0];
  _RAND_2979 = {1{`RANDOM}};
  reg_csr_2979 = _RAND_2979[31:0];
  _RAND_2980 = {1{`RANDOM}};
  reg_csr_2980 = _RAND_2980[31:0];
  _RAND_2981 = {1{`RANDOM}};
  reg_csr_2981 = _RAND_2981[31:0];
  _RAND_2982 = {1{`RANDOM}};
  reg_csr_2982 = _RAND_2982[31:0];
  _RAND_2983 = {1{`RANDOM}};
  reg_csr_2983 = _RAND_2983[31:0];
  _RAND_2984 = {1{`RANDOM}};
  reg_csr_2984 = _RAND_2984[31:0];
  _RAND_2985 = {1{`RANDOM}};
  reg_csr_2985 = _RAND_2985[31:0];
  _RAND_2986 = {1{`RANDOM}};
  reg_csr_2986 = _RAND_2986[31:0];
  _RAND_2987 = {1{`RANDOM}};
  reg_csr_2987 = _RAND_2987[31:0];
  _RAND_2988 = {1{`RANDOM}};
  reg_csr_2988 = _RAND_2988[31:0];
  _RAND_2989 = {1{`RANDOM}};
  reg_csr_2989 = _RAND_2989[31:0];
  _RAND_2990 = {1{`RANDOM}};
  reg_csr_2990 = _RAND_2990[31:0];
  _RAND_2991 = {1{`RANDOM}};
  reg_csr_2991 = _RAND_2991[31:0];
  _RAND_2992 = {1{`RANDOM}};
  reg_csr_2992 = _RAND_2992[31:0];
  _RAND_2993 = {1{`RANDOM}};
  reg_csr_2993 = _RAND_2993[31:0];
  _RAND_2994 = {1{`RANDOM}};
  reg_csr_2994 = _RAND_2994[31:0];
  _RAND_2995 = {1{`RANDOM}};
  reg_csr_2995 = _RAND_2995[31:0];
  _RAND_2996 = {1{`RANDOM}};
  reg_csr_2996 = _RAND_2996[31:0];
  _RAND_2997 = {1{`RANDOM}};
  reg_csr_2997 = _RAND_2997[31:0];
  _RAND_2998 = {1{`RANDOM}};
  reg_csr_2998 = _RAND_2998[31:0];
  _RAND_2999 = {1{`RANDOM}};
  reg_csr_2999 = _RAND_2999[31:0];
  _RAND_3000 = {1{`RANDOM}};
  reg_csr_3000 = _RAND_3000[31:0];
  _RAND_3001 = {1{`RANDOM}};
  reg_csr_3001 = _RAND_3001[31:0];
  _RAND_3002 = {1{`RANDOM}};
  reg_csr_3002 = _RAND_3002[31:0];
  _RAND_3003 = {1{`RANDOM}};
  reg_csr_3003 = _RAND_3003[31:0];
  _RAND_3004 = {1{`RANDOM}};
  reg_csr_3004 = _RAND_3004[31:0];
  _RAND_3005 = {1{`RANDOM}};
  reg_csr_3005 = _RAND_3005[31:0];
  _RAND_3006 = {1{`RANDOM}};
  reg_csr_3006 = _RAND_3006[31:0];
  _RAND_3007 = {1{`RANDOM}};
  reg_csr_3007 = _RAND_3007[31:0];
  _RAND_3008 = {1{`RANDOM}};
  reg_csr_3008 = _RAND_3008[31:0];
  _RAND_3009 = {1{`RANDOM}};
  reg_csr_3009 = _RAND_3009[31:0];
  _RAND_3010 = {1{`RANDOM}};
  reg_csr_3010 = _RAND_3010[31:0];
  _RAND_3011 = {1{`RANDOM}};
  reg_csr_3011 = _RAND_3011[31:0];
  _RAND_3012 = {1{`RANDOM}};
  reg_csr_3012 = _RAND_3012[31:0];
  _RAND_3013 = {1{`RANDOM}};
  reg_csr_3013 = _RAND_3013[31:0];
  _RAND_3014 = {1{`RANDOM}};
  reg_csr_3014 = _RAND_3014[31:0];
  _RAND_3015 = {1{`RANDOM}};
  reg_csr_3015 = _RAND_3015[31:0];
  _RAND_3016 = {1{`RANDOM}};
  reg_csr_3016 = _RAND_3016[31:0];
  _RAND_3017 = {1{`RANDOM}};
  reg_csr_3017 = _RAND_3017[31:0];
  _RAND_3018 = {1{`RANDOM}};
  reg_csr_3018 = _RAND_3018[31:0];
  _RAND_3019 = {1{`RANDOM}};
  reg_csr_3019 = _RAND_3019[31:0];
  _RAND_3020 = {1{`RANDOM}};
  reg_csr_3020 = _RAND_3020[31:0];
  _RAND_3021 = {1{`RANDOM}};
  reg_csr_3021 = _RAND_3021[31:0];
  _RAND_3022 = {1{`RANDOM}};
  reg_csr_3022 = _RAND_3022[31:0];
  _RAND_3023 = {1{`RANDOM}};
  reg_csr_3023 = _RAND_3023[31:0];
  _RAND_3024 = {1{`RANDOM}};
  reg_csr_3024 = _RAND_3024[31:0];
  _RAND_3025 = {1{`RANDOM}};
  reg_csr_3025 = _RAND_3025[31:0];
  _RAND_3026 = {1{`RANDOM}};
  reg_csr_3026 = _RAND_3026[31:0];
  _RAND_3027 = {1{`RANDOM}};
  reg_csr_3027 = _RAND_3027[31:0];
  _RAND_3028 = {1{`RANDOM}};
  reg_csr_3028 = _RAND_3028[31:0];
  _RAND_3029 = {1{`RANDOM}};
  reg_csr_3029 = _RAND_3029[31:0];
  _RAND_3030 = {1{`RANDOM}};
  reg_csr_3030 = _RAND_3030[31:0];
  _RAND_3031 = {1{`RANDOM}};
  reg_csr_3031 = _RAND_3031[31:0];
  _RAND_3032 = {1{`RANDOM}};
  reg_csr_3032 = _RAND_3032[31:0];
  _RAND_3033 = {1{`RANDOM}};
  reg_csr_3033 = _RAND_3033[31:0];
  _RAND_3034 = {1{`RANDOM}};
  reg_csr_3034 = _RAND_3034[31:0];
  _RAND_3035 = {1{`RANDOM}};
  reg_csr_3035 = _RAND_3035[31:0];
  _RAND_3036 = {1{`RANDOM}};
  reg_csr_3036 = _RAND_3036[31:0];
  _RAND_3037 = {1{`RANDOM}};
  reg_csr_3037 = _RAND_3037[31:0];
  _RAND_3038 = {1{`RANDOM}};
  reg_csr_3038 = _RAND_3038[31:0];
  _RAND_3039 = {1{`RANDOM}};
  reg_csr_3039 = _RAND_3039[31:0];
  _RAND_3040 = {1{`RANDOM}};
  reg_csr_3040 = _RAND_3040[31:0];
  _RAND_3041 = {1{`RANDOM}};
  reg_csr_3041 = _RAND_3041[31:0];
  _RAND_3042 = {1{`RANDOM}};
  reg_csr_3042 = _RAND_3042[31:0];
  _RAND_3043 = {1{`RANDOM}};
  reg_csr_3043 = _RAND_3043[31:0];
  _RAND_3044 = {1{`RANDOM}};
  reg_csr_3044 = _RAND_3044[31:0];
  _RAND_3045 = {1{`RANDOM}};
  reg_csr_3045 = _RAND_3045[31:0];
  _RAND_3046 = {1{`RANDOM}};
  reg_csr_3046 = _RAND_3046[31:0];
  _RAND_3047 = {1{`RANDOM}};
  reg_csr_3047 = _RAND_3047[31:0];
  _RAND_3048 = {1{`RANDOM}};
  reg_csr_3048 = _RAND_3048[31:0];
  _RAND_3049 = {1{`RANDOM}};
  reg_csr_3049 = _RAND_3049[31:0];
  _RAND_3050 = {1{`RANDOM}};
  reg_csr_3050 = _RAND_3050[31:0];
  _RAND_3051 = {1{`RANDOM}};
  reg_csr_3051 = _RAND_3051[31:0];
  _RAND_3052 = {1{`RANDOM}};
  reg_csr_3052 = _RAND_3052[31:0];
  _RAND_3053 = {1{`RANDOM}};
  reg_csr_3053 = _RAND_3053[31:0];
  _RAND_3054 = {1{`RANDOM}};
  reg_csr_3054 = _RAND_3054[31:0];
  _RAND_3055 = {1{`RANDOM}};
  reg_csr_3055 = _RAND_3055[31:0];
  _RAND_3056 = {1{`RANDOM}};
  reg_csr_3056 = _RAND_3056[31:0];
  _RAND_3057 = {1{`RANDOM}};
  reg_csr_3057 = _RAND_3057[31:0];
  _RAND_3058 = {1{`RANDOM}};
  reg_csr_3058 = _RAND_3058[31:0];
  _RAND_3059 = {1{`RANDOM}};
  reg_csr_3059 = _RAND_3059[31:0];
  _RAND_3060 = {1{`RANDOM}};
  reg_csr_3060 = _RAND_3060[31:0];
  _RAND_3061 = {1{`RANDOM}};
  reg_csr_3061 = _RAND_3061[31:0];
  _RAND_3062 = {1{`RANDOM}};
  reg_csr_3062 = _RAND_3062[31:0];
  _RAND_3063 = {1{`RANDOM}};
  reg_csr_3063 = _RAND_3063[31:0];
  _RAND_3064 = {1{`RANDOM}};
  reg_csr_3064 = _RAND_3064[31:0];
  _RAND_3065 = {1{`RANDOM}};
  reg_csr_3065 = _RAND_3065[31:0];
  _RAND_3066 = {1{`RANDOM}};
  reg_csr_3066 = _RAND_3066[31:0];
  _RAND_3067 = {1{`RANDOM}};
  reg_csr_3067 = _RAND_3067[31:0];
  _RAND_3068 = {1{`RANDOM}};
  reg_csr_3068 = _RAND_3068[31:0];
  _RAND_3069 = {1{`RANDOM}};
  reg_csr_3069 = _RAND_3069[31:0];
  _RAND_3070 = {1{`RANDOM}};
  reg_csr_3070 = _RAND_3070[31:0];
  _RAND_3071 = {1{`RANDOM}};
  reg_csr_3071 = _RAND_3071[31:0];
  _RAND_3072 = {1{`RANDOM}};
  reg_csr_3072 = _RAND_3072[31:0];
  _RAND_3073 = {1{`RANDOM}};
  reg_csr_3073 = _RAND_3073[31:0];
  _RAND_3074 = {1{`RANDOM}};
  reg_csr_3074 = _RAND_3074[31:0];
  _RAND_3075 = {1{`RANDOM}};
  reg_csr_3075 = _RAND_3075[31:0];
  _RAND_3076 = {1{`RANDOM}};
  reg_csr_3076 = _RAND_3076[31:0];
  _RAND_3077 = {1{`RANDOM}};
  reg_csr_3077 = _RAND_3077[31:0];
  _RAND_3078 = {1{`RANDOM}};
  reg_csr_3078 = _RAND_3078[31:0];
  _RAND_3079 = {1{`RANDOM}};
  reg_csr_3079 = _RAND_3079[31:0];
  _RAND_3080 = {1{`RANDOM}};
  reg_csr_3080 = _RAND_3080[31:0];
  _RAND_3081 = {1{`RANDOM}};
  reg_csr_3081 = _RAND_3081[31:0];
  _RAND_3082 = {1{`RANDOM}};
  reg_csr_3082 = _RAND_3082[31:0];
  _RAND_3083 = {1{`RANDOM}};
  reg_csr_3083 = _RAND_3083[31:0];
  _RAND_3084 = {1{`RANDOM}};
  reg_csr_3084 = _RAND_3084[31:0];
  _RAND_3085 = {1{`RANDOM}};
  reg_csr_3085 = _RAND_3085[31:0];
  _RAND_3086 = {1{`RANDOM}};
  reg_csr_3086 = _RAND_3086[31:0];
  _RAND_3087 = {1{`RANDOM}};
  reg_csr_3087 = _RAND_3087[31:0];
  _RAND_3088 = {1{`RANDOM}};
  reg_csr_3088 = _RAND_3088[31:0];
  _RAND_3089 = {1{`RANDOM}};
  reg_csr_3089 = _RAND_3089[31:0];
  _RAND_3090 = {1{`RANDOM}};
  reg_csr_3090 = _RAND_3090[31:0];
  _RAND_3091 = {1{`RANDOM}};
  reg_csr_3091 = _RAND_3091[31:0];
  _RAND_3092 = {1{`RANDOM}};
  reg_csr_3092 = _RAND_3092[31:0];
  _RAND_3093 = {1{`RANDOM}};
  reg_csr_3093 = _RAND_3093[31:0];
  _RAND_3094 = {1{`RANDOM}};
  reg_csr_3094 = _RAND_3094[31:0];
  _RAND_3095 = {1{`RANDOM}};
  reg_csr_3095 = _RAND_3095[31:0];
  _RAND_3096 = {1{`RANDOM}};
  reg_csr_3096 = _RAND_3096[31:0];
  _RAND_3097 = {1{`RANDOM}};
  reg_csr_3097 = _RAND_3097[31:0];
  _RAND_3098 = {1{`RANDOM}};
  reg_csr_3098 = _RAND_3098[31:0];
  _RAND_3099 = {1{`RANDOM}};
  reg_csr_3099 = _RAND_3099[31:0];
  _RAND_3100 = {1{`RANDOM}};
  reg_csr_3100 = _RAND_3100[31:0];
  _RAND_3101 = {1{`RANDOM}};
  reg_csr_3101 = _RAND_3101[31:0];
  _RAND_3102 = {1{`RANDOM}};
  reg_csr_3102 = _RAND_3102[31:0];
  _RAND_3103 = {1{`RANDOM}};
  reg_csr_3103 = _RAND_3103[31:0];
  _RAND_3104 = {1{`RANDOM}};
  reg_csr_3104 = _RAND_3104[31:0];
  _RAND_3105 = {1{`RANDOM}};
  reg_csr_3105 = _RAND_3105[31:0];
  _RAND_3106 = {1{`RANDOM}};
  reg_csr_3106 = _RAND_3106[31:0];
  _RAND_3107 = {1{`RANDOM}};
  reg_csr_3107 = _RAND_3107[31:0];
  _RAND_3108 = {1{`RANDOM}};
  reg_csr_3108 = _RAND_3108[31:0];
  _RAND_3109 = {1{`RANDOM}};
  reg_csr_3109 = _RAND_3109[31:0];
  _RAND_3110 = {1{`RANDOM}};
  reg_csr_3110 = _RAND_3110[31:0];
  _RAND_3111 = {1{`RANDOM}};
  reg_csr_3111 = _RAND_3111[31:0];
  _RAND_3112 = {1{`RANDOM}};
  reg_csr_3112 = _RAND_3112[31:0];
  _RAND_3113 = {1{`RANDOM}};
  reg_csr_3113 = _RAND_3113[31:0];
  _RAND_3114 = {1{`RANDOM}};
  reg_csr_3114 = _RAND_3114[31:0];
  _RAND_3115 = {1{`RANDOM}};
  reg_csr_3115 = _RAND_3115[31:0];
  _RAND_3116 = {1{`RANDOM}};
  reg_csr_3116 = _RAND_3116[31:0];
  _RAND_3117 = {1{`RANDOM}};
  reg_csr_3117 = _RAND_3117[31:0];
  _RAND_3118 = {1{`RANDOM}};
  reg_csr_3118 = _RAND_3118[31:0];
  _RAND_3119 = {1{`RANDOM}};
  reg_csr_3119 = _RAND_3119[31:0];
  _RAND_3120 = {1{`RANDOM}};
  reg_csr_3120 = _RAND_3120[31:0];
  _RAND_3121 = {1{`RANDOM}};
  reg_csr_3121 = _RAND_3121[31:0];
  _RAND_3122 = {1{`RANDOM}};
  reg_csr_3122 = _RAND_3122[31:0];
  _RAND_3123 = {1{`RANDOM}};
  reg_csr_3123 = _RAND_3123[31:0];
  _RAND_3124 = {1{`RANDOM}};
  reg_csr_3124 = _RAND_3124[31:0];
  _RAND_3125 = {1{`RANDOM}};
  reg_csr_3125 = _RAND_3125[31:0];
  _RAND_3126 = {1{`RANDOM}};
  reg_csr_3126 = _RAND_3126[31:0];
  _RAND_3127 = {1{`RANDOM}};
  reg_csr_3127 = _RAND_3127[31:0];
  _RAND_3128 = {1{`RANDOM}};
  reg_csr_3128 = _RAND_3128[31:0];
  _RAND_3129 = {1{`RANDOM}};
  reg_csr_3129 = _RAND_3129[31:0];
  _RAND_3130 = {1{`RANDOM}};
  reg_csr_3130 = _RAND_3130[31:0];
  _RAND_3131 = {1{`RANDOM}};
  reg_csr_3131 = _RAND_3131[31:0];
  _RAND_3132 = {1{`RANDOM}};
  reg_csr_3132 = _RAND_3132[31:0];
  _RAND_3133 = {1{`RANDOM}};
  reg_csr_3133 = _RAND_3133[31:0];
  _RAND_3134 = {1{`RANDOM}};
  reg_csr_3134 = _RAND_3134[31:0];
  _RAND_3135 = {1{`RANDOM}};
  reg_csr_3135 = _RAND_3135[31:0];
  _RAND_3136 = {1{`RANDOM}};
  reg_csr_3136 = _RAND_3136[31:0];
  _RAND_3137 = {1{`RANDOM}};
  reg_csr_3137 = _RAND_3137[31:0];
  _RAND_3138 = {1{`RANDOM}};
  reg_csr_3138 = _RAND_3138[31:0];
  _RAND_3139 = {1{`RANDOM}};
  reg_csr_3139 = _RAND_3139[31:0];
  _RAND_3140 = {1{`RANDOM}};
  reg_csr_3140 = _RAND_3140[31:0];
  _RAND_3141 = {1{`RANDOM}};
  reg_csr_3141 = _RAND_3141[31:0];
  _RAND_3142 = {1{`RANDOM}};
  reg_csr_3142 = _RAND_3142[31:0];
  _RAND_3143 = {1{`RANDOM}};
  reg_csr_3143 = _RAND_3143[31:0];
  _RAND_3144 = {1{`RANDOM}};
  reg_csr_3144 = _RAND_3144[31:0];
  _RAND_3145 = {1{`RANDOM}};
  reg_csr_3145 = _RAND_3145[31:0];
  _RAND_3146 = {1{`RANDOM}};
  reg_csr_3146 = _RAND_3146[31:0];
  _RAND_3147 = {1{`RANDOM}};
  reg_csr_3147 = _RAND_3147[31:0];
  _RAND_3148 = {1{`RANDOM}};
  reg_csr_3148 = _RAND_3148[31:0];
  _RAND_3149 = {1{`RANDOM}};
  reg_csr_3149 = _RAND_3149[31:0];
  _RAND_3150 = {1{`RANDOM}};
  reg_csr_3150 = _RAND_3150[31:0];
  _RAND_3151 = {1{`RANDOM}};
  reg_csr_3151 = _RAND_3151[31:0];
  _RAND_3152 = {1{`RANDOM}};
  reg_csr_3152 = _RAND_3152[31:0];
  _RAND_3153 = {1{`RANDOM}};
  reg_csr_3153 = _RAND_3153[31:0];
  _RAND_3154 = {1{`RANDOM}};
  reg_csr_3154 = _RAND_3154[31:0];
  _RAND_3155 = {1{`RANDOM}};
  reg_csr_3155 = _RAND_3155[31:0];
  _RAND_3156 = {1{`RANDOM}};
  reg_csr_3156 = _RAND_3156[31:0];
  _RAND_3157 = {1{`RANDOM}};
  reg_csr_3157 = _RAND_3157[31:0];
  _RAND_3158 = {1{`RANDOM}};
  reg_csr_3158 = _RAND_3158[31:0];
  _RAND_3159 = {1{`RANDOM}};
  reg_csr_3159 = _RAND_3159[31:0];
  _RAND_3160 = {1{`RANDOM}};
  reg_csr_3160 = _RAND_3160[31:0];
  _RAND_3161 = {1{`RANDOM}};
  reg_csr_3161 = _RAND_3161[31:0];
  _RAND_3162 = {1{`RANDOM}};
  reg_csr_3162 = _RAND_3162[31:0];
  _RAND_3163 = {1{`RANDOM}};
  reg_csr_3163 = _RAND_3163[31:0];
  _RAND_3164 = {1{`RANDOM}};
  reg_csr_3164 = _RAND_3164[31:0];
  _RAND_3165 = {1{`RANDOM}};
  reg_csr_3165 = _RAND_3165[31:0];
  _RAND_3166 = {1{`RANDOM}};
  reg_csr_3166 = _RAND_3166[31:0];
  _RAND_3167 = {1{`RANDOM}};
  reg_csr_3167 = _RAND_3167[31:0];
  _RAND_3168 = {1{`RANDOM}};
  reg_csr_3168 = _RAND_3168[31:0];
  _RAND_3169 = {1{`RANDOM}};
  reg_csr_3169 = _RAND_3169[31:0];
  _RAND_3170 = {1{`RANDOM}};
  reg_csr_3170 = _RAND_3170[31:0];
  _RAND_3171 = {1{`RANDOM}};
  reg_csr_3171 = _RAND_3171[31:0];
  _RAND_3172 = {1{`RANDOM}};
  reg_csr_3172 = _RAND_3172[31:0];
  _RAND_3173 = {1{`RANDOM}};
  reg_csr_3173 = _RAND_3173[31:0];
  _RAND_3174 = {1{`RANDOM}};
  reg_csr_3174 = _RAND_3174[31:0];
  _RAND_3175 = {1{`RANDOM}};
  reg_csr_3175 = _RAND_3175[31:0];
  _RAND_3176 = {1{`RANDOM}};
  reg_csr_3176 = _RAND_3176[31:0];
  _RAND_3177 = {1{`RANDOM}};
  reg_csr_3177 = _RAND_3177[31:0];
  _RAND_3178 = {1{`RANDOM}};
  reg_csr_3178 = _RAND_3178[31:0];
  _RAND_3179 = {1{`RANDOM}};
  reg_csr_3179 = _RAND_3179[31:0];
  _RAND_3180 = {1{`RANDOM}};
  reg_csr_3180 = _RAND_3180[31:0];
  _RAND_3181 = {1{`RANDOM}};
  reg_csr_3181 = _RAND_3181[31:0];
  _RAND_3182 = {1{`RANDOM}};
  reg_csr_3182 = _RAND_3182[31:0];
  _RAND_3183 = {1{`RANDOM}};
  reg_csr_3183 = _RAND_3183[31:0];
  _RAND_3184 = {1{`RANDOM}};
  reg_csr_3184 = _RAND_3184[31:0];
  _RAND_3185 = {1{`RANDOM}};
  reg_csr_3185 = _RAND_3185[31:0];
  _RAND_3186 = {1{`RANDOM}};
  reg_csr_3186 = _RAND_3186[31:0];
  _RAND_3187 = {1{`RANDOM}};
  reg_csr_3187 = _RAND_3187[31:0];
  _RAND_3188 = {1{`RANDOM}};
  reg_csr_3188 = _RAND_3188[31:0];
  _RAND_3189 = {1{`RANDOM}};
  reg_csr_3189 = _RAND_3189[31:0];
  _RAND_3190 = {1{`RANDOM}};
  reg_csr_3190 = _RAND_3190[31:0];
  _RAND_3191 = {1{`RANDOM}};
  reg_csr_3191 = _RAND_3191[31:0];
  _RAND_3192 = {1{`RANDOM}};
  reg_csr_3192 = _RAND_3192[31:0];
  _RAND_3193 = {1{`RANDOM}};
  reg_csr_3193 = _RAND_3193[31:0];
  _RAND_3194 = {1{`RANDOM}};
  reg_csr_3194 = _RAND_3194[31:0];
  _RAND_3195 = {1{`RANDOM}};
  reg_csr_3195 = _RAND_3195[31:0];
  _RAND_3196 = {1{`RANDOM}};
  reg_csr_3196 = _RAND_3196[31:0];
  _RAND_3197 = {1{`RANDOM}};
  reg_csr_3197 = _RAND_3197[31:0];
  _RAND_3198 = {1{`RANDOM}};
  reg_csr_3198 = _RAND_3198[31:0];
  _RAND_3199 = {1{`RANDOM}};
  reg_csr_3199 = _RAND_3199[31:0];
  _RAND_3200 = {1{`RANDOM}};
  reg_csr_3200 = _RAND_3200[31:0];
  _RAND_3201 = {1{`RANDOM}};
  reg_csr_3201 = _RAND_3201[31:0];
  _RAND_3202 = {1{`RANDOM}};
  reg_csr_3202 = _RAND_3202[31:0];
  _RAND_3203 = {1{`RANDOM}};
  reg_csr_3203 = _RAND_3203[31:0];
  _RAND_3204 = {1{`RANDOM}};
  reg_csr_3204 = _RAND_3204[31:0];
  _RAND_3205 = {1{`RANDOM}};
  reg_csr_3205 = _RAND_3205[31:0];
  _RAND_3206 = {1{`RANDOM}};
  reg_csr_3206 = _RAND_3206[31:0];
  _RAND_3207 = {1{`RANDOM}};
  reg_csr_3207 = _RAND_3207[31:0];
  _RAND_3208 = {1{`RANDOM}};
  reg_csr_3208 = _RAND_3208[31:0];
  _RAND_3209 = {1{`RANDOM}};
  reg_csr_3209 = _RAND_3209[31:0];
  _RAND_3210 = {1{`RANDOM}};
  reg_csr_3210 = _RAND_3210[31:0];
  _RAND_3211 = {1{`RANDOM}};
  reg_csr_3211 = _RAND_3211[31:0];
  _RAND_3212 = {1{`RANDOM}};
  reg_csr_3212 = _RAND_3212[31:0];
  _RAND_3213 = {1{`RANDOM}};
  reg_csr_3213 = _RAND_3213[31:0];
  _RAND_3214 = {1{`RANDOM}};
  reg_csr_3214 = _RAND_3214[31:0];
  _RAND_3215 = {1{`RANDOM}};
  reg_csr_3215 = _RAND_3215[31:0];
  _RAND_3216 = {1{`RANDOM}};
  reg_csr_3216 = _RAND_3216[31:0];
  _RAND_3217 = {1{`RANDOM}};
  reg_csr_3217 = _RAND_3217[31:0];
  _RAND_3218 = {1{`RANDOM}};
  reg_csr_3218 = _RAND_3218[31:0];
  _RAND_3219 = {1{`RANDOM}};
  reg_csr_3219 = _RAND_3219[31:0];
  _RAND_3220 = {1{`RANDOM}};
  reg_csr_3220 = _RAND_3220[31:0];
  _RAND_3221 = {1{`RANDOM}};
  reg_csr_3221 = _RAND_3221[31:0];
  _RAND_3222 = {1{`RANDOM}};
  reg_csr_3222 = _RAND_3222[31:0];
  _RAND_3223 = {1{`RANDOM}};
  reg_csr_3223 = _RAND_3223[31:0];
  _RAND_3224 = {1{`RANDOM}};
  reg_csr_3224 = _RAND_3224[31:0];
  _RAND_3225 = {1{`RANDOM}};
  reg_csr_3225 = _RAND_3225[31:0];
  _RAND_3226 = {1{`RANDOM}};
  reg_csr_3226 = _RAND_3226[31:0];
  _RAND_3227 = {1{`RANDOM}};
  reg_csr_3227 = _RAND_3227[31:0];
  _RAND_3228 = {1{`RANDOM}};
  reg_csr_3228 = _RAND_3228[31:0];
  _RAND_3229 = {1{`RANDOM}};
  reg_csr_3229 = _RAND_3229[31:0];
  _RAND_3230 = {1{`RANDOM}};
  reg_csr_3230 = _RAND_3230[31:0];
  _RAND_3231 = {1{`RANDOM}};
  reg_csr_3231 = _RAND_3231[31:0];
  _RAND_3232 = {1{`RANDOM}};
  reg_csr_3232 = _RAND_3232[31:0];
  _RAND_3233 = {1{`RANDOM}};
  reg_csr_3233 = _RAND_3233[31:0];
  _RAND_3234 = {1{`RANDOM}};
  reg_csr_3234 = _RAND_3234[31:0];
  _RAND_3235 = {1{`RANDOM}};
  reg_csr_3235 = _RAND_3235[31:0];
  _RAND_3236 = {1{`RANDOM}};
  reg_csr_3236 = _RAND_3236[31:0];
  _RAND_3237 = {1{`RANDOM}};
  reg_csr_3237 = _RAND_3237[31:0];
  _RAND_3238 = {1{`RANDOM}};
  reg_csr_3238 = _RAND_3238[31:0];
  _RAND_3239 = {1{`RANDOM}};
  reg_csr_3239 = _RAND_3239[31:0];
  _RAND_3240 = {1{`RANDOM}};
  reg_csr_3240 = _RAND_3240[31:0];
  _RAND_3241 = {1{`RANDOM}};
  reg_csr_3241 = _RAND_3241[31:0];
  _RAND_3242 = {1{`RANDOM}};
  reg_csr_3242 = _RAND_3242[31:0];
  _RAND_3243 = {1{`RANDOM}};
  reg_csr_3243 = _RAND_3243[31:0];
  _RAND_3244 = {1{`RANDOM}};
  reg_csr_3244 = _RAND_3244[31:0];
  _RAND_3245 = {1{`RANDOM}};
  reg_csr_3245 = _RAND_3245[31:0];
  _RAND_3246 = {1{`RANDOM}};
  reg_csr_3246 = _RAND_3246[31:0];
  _RAND_3247 = {1{`RANDOM}};
  reg_csr_3247 = _RAND_3247[31:0];
  _RAND_3248 = {1{`RANDOM}};
  reg_csr_3248 = _RAND_3248[31:0];
  _RAND_3249 = {1{`RANDOM}};
  reg_csr_3249 = _RAND_3249[31:0];
  _RAND_3250 = {1{`RANDOM}};
  reg_csr_3250 = _RAND_3250[31:0];
  _RAND_3251 = {1{`RANDOM}};
  reg_csr_3251 = _RAND_3251[31:0];
  _RAND_3252 = {1{`RANDOM}};
  reg_csr_3252 = _RAND_3252[31:0];
  _RAND_3253 = {1{`RANDOM}};
  reg_csr_3253 = _RAND_3253[31:0];
  _RAND_3254 = {1{`RANDOM}};
  reg_csr_3254 = _RAND_3254[31:0];
  _RAND_3255 = {1{`RANDOM}};
  reg_csr_3255 = _RAND_3255[31:0];
  _RAND_3256 = {1{`RANDOM}};
  reg_csr_3256 = _RAND_3256[31:0];
  _RAND_3257 = {1{`RANDOM}};
  reg_csr_3257 = _RAND_3257[31:0];
  _RAND_3258 = {1{`RANDOM}};
  reg_csr_3258 = _RAND_3258[31:0];
  _RAND_3259 = {1{`RANDOM}};
  reg_csr_3259 = _RAND_3259[31:0];
  _RAND_3260 = {1{`RANDOM}};
  reg_csr_3260 = _RAND_3260[31:0];
  _RAND_3261 = {1{`RANDOM}};
  reg_csr_3261 = _RAND_3261[31:0];
  _RAND_3262 = {1{`RANDOM}};
  reg_csr_3262 = _RAND_3262[31:0];
  _RAND_3263 = {1{`RANDOM}};
  reg_csr_3263 = _RAND_3263[31:0];
  _RAND_3264 = {1{`RANDOM}};
  reg_csr_3264 = _RAND_3264[31:0];
  _RAND_3265 = {1{`RANDOM}};
  reg_csr_3265 = _RAND_3265[31:0];
  _RAND_3266 = {1{`RANDOM}};
  reg_csr_3266 = _RAND_3266[31:0];
  _RAND_3267 = {1{`RANDOM}};
  reg_csr_3267 = _RAND_3267[31:0];
  _RAND_3268 = {1{`RANDOM}};
  reg_csr_3268 = _RAND_3268[31:0];
  _RAND_3269 = {1{`RANDOM}};
  reg_csr_3269 = _RAND_3269[31:0];
  _RAND_3270 = {1{`RANDOM}};
  reg_csr_3270 = _RAND_3270[31:0];
  _RAND_3271 = {1{`RANDOM}};
  reg_csr_3271 = _RAND_3271[31:0];
  _RAND_3272 = {1{`RANDOM}};
  reg_csr_3272 = _RAND_3272[31:0];
  _RAND_3273 = {1{`RANDOM}};
  reg_csr_3273 = _RAND_3273[31:0];
  _RAND_3274 = {1{`RANDOM}};
  reg_csr_3274 = _RAND_3274[31:0];
  _RAND_3275 = {1{`RANDOM}};
  reg_csr_3275 = _RAND_3275[31:0];
  _RAND_3276 = {1{`RANDOM}};
  reg_csr_3276 = _RAND_3276[31:0];
  _RAND_3277 = {1{`RANDOM}};
  reg_csr_3277 = _RAND_3277[31:0];
  _RAND_3278 = {1{`RANDOM}};
  reg_csr_3278 = _RAND_3278[31:0];
  _RAND_3279 = {1{`RANDOM}};
  reg_csr_3279 = _RAND_3279[31:0];
  _RAND_3280 = {1{`RANDOM}};
  reg_csr_3280 = _RAND_3280[31:0];
  _RAND_3281 = {1{`RANDOM}};
  reg_csr_3281 = _RAND_3281[31:0];
  _RAND_3282 = {1{`RANDOM}};
  reg_csr_3282 = _RAND_3282[31:0];
  _RAND_3283 = {1{`RANDOM}};
  reg_csr_3283 = _RAND_3283[31:0];
  _RAND_3284 = {1{`RANDOM}};
  reg_csr_3284 = _RAND_3284[31:0];
  _RAND_3285 = {1{`RANDOM}};
  reg_csr_3285 = _RAND_3285[31:0];
  _RAND_3286 = {1{`RANDOM}};
  reg_csr_3286 = _RAND_3286[31:0];
  _RAND_3287 = {1{`RANDOM}};
  reg_csr_3287 = _RAND_3287[31:0];
  _RAND_3288 = {1{`RANDOM}};
  reg_csr_3288 = _RAND_3288[31:0];
  _RAND_3289 = {1{`RANDOM}};
  reg_csr_3289 = _RAND_3289[31:0];
  _RAND_3290 = {1{`RANDOM}};
  reg_csr_3290 = _RAND_3290[31:0];
  _RAND_3291 = {1{`RANDOM}};
  reg_csr_3291 = _RAND_3291[31:0];
  _RAND_3292 = {1{`RANDOM}};
  reg_csr_3292 = _RAND_3292[31:0];
  _RAND_3293 = {1{`RANDOM}};
  reg_csr_3293 = _RAND_3293[31:0];
  _RAND_3294 = {1{`RANDOM}};
  reg_csr_3294 = _RAND_3294[31:0];
  _RAND_3295 = {1{`RANDOM}};
  reg_csr_3295 = _RAND_3295[31:0];
  _RAND_3296 = {1{`RANDOM}};
  reg_csr_3296 = _RAND_3296[31:0];
  _RAND_3297 = {1{`RANDOM}};
  reg_csr_3297 = _RAND_3297[31:0];
  _RAND_3298 = {1{`RANDOM}};
  reg_csr_3298 = _RAND_3298[31:0];
  _RAND_3299 = {1{`RANDOM}};
  reg_csr_3299 = _RAND_3299[31:0];
  _RAND_3300 = {1{`RANDOM}};
  reg_csr_3300 = _RAND_3300[31:0];
  _RAND_3301 = {1{`RANDOM}};
  reg_csr_3301 = _RAND_3301[31:0];
  _RAND_3302 = {1{`RANDOM}};
  reg_csr_3302 = _RAND_3302[31:0];
  _RAND_3303 = {1{`RANDOM}};
  reg_csr_3303 = _RAND_3303[31:0];
  _RAND_3304 = {1{`RANDOM}};
  reg_csr_3304 = _RAND_3304[31:0];
  _RAND_3305 = {1{`RANDOM}};
  reg_csr_3305 = _RAND_3305[31:0];
  _RAND_3306 = {1{`RANDOM}};
  reg_csr_3306 = _RAND_3306[31:0];
  _RAND_3307 = {1{`RANDOM}};
  reg_csr_3307 = _RAND_3307[31:0];
  _RAND_3308 = {1{`RANDOM}};
  reg_csr_3308 = _RAND_3308[31:0];
  _RAND_3309 = {1{`RANDOM}};
  reg_csr_3309 = _RAND_3309[31:0];
  _RAND_3310 = {1{`RANDOM}};
  reg_csr_3310 = _RAND_3310[31:0];
  _RAND_3311 = {1{`RANDOM}};
  reg_csr_3311 = _RAND_3311[31:0];
  _RAND_3312 = {1{`RANDOM}};
  reg_csr_3312 = _RAND_3312[31:0];
  _RAND_3313 = {1{`RANDOM}};
  reg_csr_3313 = _RAND_3313[31:0];
  _RAND_3314 = {1{`RANDOM}};
  reg_csr_3314 = _RAND_3314[31:0];
  _RAND_3315 = {1{`RANDOM}};
  reg_csr_3315 = _RAND_3315[31:0];
  _RAND_3316 = {1{`RANDOM}};
  reg_csr_3316 = _RAND_3316[31:0];
  _RAND_3317 = {1{`RANDOM}};
  reg_csr_3317 = _RAND_3317[31:0];
  _RAND_3318 = {1{`RANDOM}};
  reg_csr_3318 = _RAND_3318[31:0];
  _RAND_3319 = {1{`RANDOM}};
  reg_csr_3319 = _RAND_3319[31:0];
  _RAND_3320 = {1{`RANDOM}};
  reg_csr_3320 = _RAND_3320[31:0];
  _RAND_3321 = {1{`RANDOM}};
  reg_csr_3321 = _RAND_3321[31:0];
  _RAND_3322 = {1{`RANDOM}};
  reg_csr_3322 = _RAND_3322[31:0];
  _RAND_3323 = {1{`RANDOM}};
  reg_csr_3323 = _RAND_3323[31:0];
  _RAND_3324 = {1{`RANDOM}};
  reg_csr_3324 = _RAND_3324[31:0];
  _RAND_3325 = {1{`RANDOM}};
  reg_csr_3325 = _RAND_3325[31:0];
  _RAND_3326 = {1{`RANDOM}};
  reg_csr_3326 = _RAND_3326[31:0];
  _RAND_3327 = {1{`RANDOM}};
  reg_csr_3327 = _RAND_3327[31:0];
  _RAND_3328 = {1{`RANDOM}};
  reg_csr_3328 = _RAND_3328[31:0];
  _RAND_3329 = {1{`RANDOM}};
  reg_csr_3329 = _RAND_3329[31:0];
  _RAND_3330 = {1{`RANDOM}};
  reg_csr_3330 = _RAND_3330[31:0];
  _RAND_3331 = {1{`RANDOM}};
  reg_csr_3331 = _RAND_3331[31:0];
  _RAND_3332 = {1{`RANDOM}};
  reg_csr_3332 = _RAND_3332[31:0];
  _RAND_3333 = {1{`RANDOM}};
  reg_csr_3333 = _RAND_3333[31:0];
  _RAND_3334 = {1{`RANDOM}};
  reg_csr_3334 = _RAND_3334[31:0];
  _RAND_3335 = {1{`RANDOM}};
  reg_csr_3335 = _RAND_3335[31:0];
  _RAND_3336 = {1{`RANDOM}};
  reg_csr_3336 = _RAND_3336[31:0];
  _RAND_3337 = {1{`RANDOM}};
  reg_csr_3337 = _RAND_3337[31:0];
  _RAND_3338 = {1{`RANDOM}};
  reg_csr_3338 = _RAND_3338[31:0];
  _RAND_3339 = {1{`RANDOM}};
  reg_csr_3339 = _RAND_3339[31:0];
  _RAND_3340 = {1{`RANDOM}};
  reg_csr_3340 = _RAND_3340[31:0];
  _RAND_3341 = {1{`RANDOM}};
  reg_csr_3341 = _RAND_3341[31:0];
  _RAND_3342 = {1{`RANDOM}};
  reg_csr_3342 = _RAND_3342[31:0];
  _RAND_3343 = {1{`RANDOM}};
  reg_csr_3343 = _RAND_3343[31:0];
  _RAND_3344 = {1{`RANDOM}};
  reg_csr_3344 = _RAND_3344[31:0];
  _RAND_3345 = {1{`RANDOM}};
  reg_csr_3345 = _RAND_3345[31:0];
  _RAND_3346 = {1{`RANDOM}};
  reg_csr_3346 = _RAND_3346[31:0];
  _RAND_3347 = {1{`RANDOM}};
  reg_csr_3347 = _RAND_3347[31:0];
  _RAND_3348 = {1{`RANDOM}};
  reg_csr_3348 = _RAND_3348[31:0];
  _RAND_3349 = {1{`RANDOM}};
  reg_csr_3349 = _RAND_3349[31:0];
  _RAND_3350 = {1{`RANDOM}};
  reg_csr_3350 = _RAND_3350[31:0];
  _RAND_3351 = {1{`RANDOM}};
  reg_csr_3351 = _RAND_3351[31:0];
  _RAND_3352 = {1{`RANDOM}};
  reg_csr_3352 = _RAND_3352[31:0];
  _RAND_3353 = {1{`RANDOM}};
  reg_csr_3353 = _RAND_3353[31:0];
  _RAND_3354 = {1{`RANDOM}};
  reg_csr_3354 = _RAND_3354[31:0];
  _RAND_3355 = {1{`RANDOM}};
  reg_csr_3355 = _RAND_3355[31:0];
  _RAND_3356 = {1{`RANDOM}};
  reg_csr_3356 = _RAND_3356[31:0];
  _RAND_3357 = {1{`RANDOM}};
  reg_csr_3357 = _RAND_3357[31:0];
  _RAND_3358 = {1{`RANDOM}};
  reg_csr_3358 = _RAND_3358[31:0];
  _RAND_3359 = {1{`RANDOM}};
  reg_csr_3359 = _RAND_3359[31:0];
  _RAND_3360 = {1{`RANDOM}};
  reg_csr_3360 = _RAND_3360[31:0];
  _RAND_3361 = {1{`RANDOM}};
  reg_csr_3361 = _RAND_3361[31:0];
  _RAND_3362 = {1{`RANDOM}};
  reg_csr_3362 = _RAND_3362[31:0];
  _RAND_3363 = {1{`RANDOM}};
  reg_csr_3363 = _RAND_3363[31:0];
  _RAND_3364 = {1{`RANDOM}};
  reg_csr_3364 = _RAND_3364[31:0];
  _RAND_3365 = {1{`RANDOM}};
  reg_csr_3365 = _RAND_3365[31:0];
  _RAND_3366 = {1{`RANDOM}};
  reg_csr_3366 = _RAND_3366[31:0];
  _RAND_3367 = {1{`RANDOM}};
  reg_csr_3367 = _RAND_3367[31:0];
  _RAND_3368 = {1{`RANDOM}};
  reg_csr_3368 = _RAND_3368[31:0];
  _RAND_3369 = {1{`RANDOM}};
  reg_csr_3369 = _RAND_3369[31:0];
  _RAND_3370 = {1{`RANDOM}};
  reg_csr_3370 = _RAND_3370[31:0];
  _RAND_3371 = {1{`RANDOM}};
  reg_csr_3371 = _RAND_3371[31:0];
  _RAND_3372 = {1{`RANDOM}};
  reg_csr_3372 = _RAND_3372[31:0];
  _RAND_3373 = {1{`RANDOM}};
  reg_csr_3373 = _RAND_3373[31:0];
  _RAND_3374 = {1{`RANDOM}};
  reg_csr_3374 = _RAND_3374[31:0];
  _RAND_3375 = {1{`RANDOM}};
  reg_csr_3375 = _RAND_3375[31:0];
  _RAND_3376 = {1{`RANDOM}};
  reg_csr_3376 = _RAND_3376[31:0];
  _RAND_3377 = {1{`RANDOM}};
  reg_csr_3377 = _RAND_3377[31:0];
  _RAND_3378 = {1{`RANDOM}};
  reg_csr_3378 = _RAND_3378[31:0];
  _RAND_3379 = {1{`RANDOM}};
  reg_csr_3379 = _RAND_3379[31:0];
  _RAND_3380 = {1{`RANDOM}};
  reg_csr_3380 = _RAND_3380[31:0];
  _RAND_3381 = {1{`RANDOM}};
  reg_csr_3381 = _RAND_3381[31:0];
  _RAND_3382 = {1{`RANDOM}};
  reg_csr_3382 = _RAND_3382[31:0];
  _RAND_3383 = {1{`RANDOM}};
  reg_csr_3383 = _RAND_3383[31:0];
  _RAND_3384 = {1{`RANDOM}};
  reg_csr_3384 = _RAND_3384[31:0];
  _RAND_3385 = {1{`RANDOM}};
  reg_csr_3385 = _RAND_3385[31:0];
  _RAND_3386 = {1{`RANDOM}};
  reg_csr_3386 = _RAND_3386[31:0];
  _RAND_3387 = {1{`RANDOM}};
  reg_csr_3387 = _RAND_3387[31:0];
  _RAND_3388 = {1{`RANDOM}};
  reg_csr_3388 = _RAND_3388[31:0];
  _RAND_3389 = {1{`RANDOM}};
  reg_csr_3389 = _RAND_3389[31:0];
  _RAND_3390 = {1{`RANDOM}};
  reg_csr_3390 = _RAND_3390[31:0];
  _RAND_3391 = {1{`RANDOM}};
  reg_csr_3391 = _RAND_3391[31:0];
  _RAND_3392 = {1{`RANDOM}};
  reg_csr_3392 = _RAND_3392[31:0];
  _RAND_3393 = {1{`RANDOM}};
  reg_csr_3393 = _RAND_3393[31:0];
  _RAND_3394 = {1{`RANDOM}};
  reg_csr_3394 = _RAND_3394[31:0];
  _RAND_3395 = {1{`RANDOM}};
  reg_csr_3395 = _RAND_3395[31:0];
  _RAND_3396 = {1{`RANDOM}};
  reg_csr_3396 = _RAND_3396[31:0];
  _RAND_3397 = {1{`RANDOM}};
  reg_csr_3397 = _RAND_3397[31:0];
  _RAND_3398 = {1{`RANDOM}};
  reg_csr_3398 = _RAND_3398[31:0];
  _RAND_3399 = {1{`RANDOM}};
  reg_csr_3399 = _RAND_3399[31:0];
  _RAND_3400 = {1{`RANDOM}};
  reg_csr_3400 = _RAND_3400[31:0];
  _RAND_3401 = {1{`RANDOM}};
  reg_csr_3401 = _RAND_3401[31:0];
  _RAND_3402 = {1{`RANDOM}};
  reg_csr_3402 = _RAND_3402[31:0];
  _RAND_3403 = {1{`RANDOM}};
  reg_csr_3403 = _RAND_3403[31:0];
  _RAND_3404 = {1{`RANDOM}};
  reg_csr_3404 = _RAND_3404[31:0];
  _RAND_3405 = {1{`RANDOM}};
  reg_csr_3405 = _RAND_3405[31:0];
  _RAND_3406 = {1{`RANDOM}};
  reg_csr_3406 = _RAND_3406[31:0];
  _RAND_3407 = {1{`RANDOM}};
  reg_csr_3407 = _RAND_3407[31:0];
  _RAND_3408 = {1{`RANDOM}};
  reg_csr_3408 = _RAND_3408[31:0];
  _RAND_3409 = {1{`RANDOM}};
  reg_csr_3409 = _RAND_3409[31:0];
  _RAND_3410 = {1{`RANDOM}};
  reg_csr_3410 = _RAND_3410[31:0];
  _RAND_3411 = {1{`RANDOM}};
  reg_csr_3411 = _RAND_3411[31:0];
  _RAND_3412 = {1{`RANDOM}};
  reg_csr_3412 = _RAND_3412[31:0];
  _RAND_3413 = {1{`RANDOM}};
  reg_csr_3413 = _RAND_3413[31:0];
  _RAND_3414 = {1{`RANDOM}};
  reg_csr_3414 = _RAND_3414[31:0];
  _RAND_3415 = {1{`RANDOM}};
  reg_csr_3415 = _RAND_3415[31:0];
  _RAND_3416 = {1{`RANDOM}};
  reg_csr_3416 = _RAND_3416[31:0];
  _RAND_3417 = {1{`RANDOM}};
  reg_csr_3417 = _RAND_3417[31:0];
  _RAND_3418 = {1{`RANDOM}};
  reg_csr_3418 = _RAND_3418[31:0];
  _RAND_3419 = {1{`RANDOM}};
  reg_csr_3419 = _RAND_3419[31:0];
  _RAND_3420 = {1{`RANDOM}};
  reg_csr_3420 = _RAND_3420[31:0];
  _RAND_3421 = {1{`RANDOM}};
  reg_csr_3421 = _RAND_3421[31:0];
  _RAND_3422 = {1{`RANDOM}};
  reg_csr_3422 = _RAND_3422[31:0];
  _RAND_3423 = {1{`RANDOM}};
  reg_csr_3423 = _RAND_3423[31:0];
  _RAND_3424 = {1{`RANDOM}};
  reg_csr_3424 = _RAND_3424[31:0];
  _RAND_3425 = {1{`RANDOM}};
  reg_csr_3425 = _RAND_3425[31:0];
  _RAND_3426 = {1{`RANDOM}};
  reg_csr_3426 = _RAND_3426[31:0];
  _RAND_3427 = {1{`RANDOM}};
  reg_csr_3427 = _RAND_3427[31:0];
  _RAND_3428 = {1{`RANDOM}};
  reg_csr_3428 = _RAND_3428[31:0];
  _RAND_3429 = {1{`RANDOM}};
  reg_csr_3429 = _RAND_3429[31:0];
  _RAND_3430 = {1{`RANDOM}};
  reg_csr_3430 = _RAND_3430[31:0];
  _RAND_3431 = {1{`RANDOM}};
  reg_csr_3431 = _RAND_3431[31:0];
  _RAND_3432 = {1{`RANDOM}};
  reg_csr_3432 = _RAND_3432[31:0];
  _RAND_3433 = {1{`RANDOM}};
  reg_csr_3433 = _RAND_3433[31:0];
  _RAND_3434 = {1{`RANDOM}};
  reg_csr_3434 = _RAND_3434[31:0];
  _RAND_3435 = {1{`RANDOM}};
  reg_csr_3435 = _RAND_3435[31:0];
  _RAND_3436 = {1{`RANDOM}};
  reg_csr_3436 = _RAND_3436[31:0];
  _RAND_3437 = {1{`RANDOM}};
  reg_csr_3437 = _RAND_3437[31:0];
  _RAND_3438 = {1{`RANDOM}};
  reg_csr_3438 = _RAND_3438[31:0];
  _RAND_3439 = {1{`RANDOM}};
  reg_csr_3439 = _RAND_3439[31:0];
  _RAND_3440 = {1{`RANDOM}};
  reg_csr_3440 = _RAND_3440[31:0];
  _RAND_3441 = {1{`RANDOM}};
  reg_csr_3441 = _RAND_3441[31:0];
  _RAND_3442 = {1{`RANDOM}};
  reg_csr_3442 = _RAND_3442[31:0];
  _RAND_3443 = {1{`RANDOM}};
  reg_csr_3443 = _RAND_3443[31:0];
  _RAND_3444 = {1{`RANDOM}};
  reg_csr_3444 = _RAND_3444[31:0];
  _RAND_3445 = {1{`RANDOM}};
  reg_csr_3445 = _RAND_3445[31:0];
  _RAND_3446 = {1{`RANDOM}};
  reg_csr_3446 = _RAND_3446[31:0];
  _RAND_3447 = {1{`RANDOM}};
  reg_csr_3447 = _RAND_3447[31:0];
  _RAND_3448 = {1{`RANDOM}};
  reg_csr_3448 = _RAND_3448[31:0];
  _RAND_3449 = {1{`RANDOM}};
  reg_csr_3449 = _RAND_3449[31:0];
  _RAND_3450 = {1{`RANDOM}};
  reg_csr_3450 = _RAND_3450[31:0];
  _RAND_3451 = {1{`RANDOM}};
  reg_csr_3451 = _RAND_3451[31:0];
  _RAND_3452 = {1{`RANDOM}};
  reg_csr_3452 = _RAND_3452[31:0];
  _RAND_3453 = {1{`RANDOM}};
  reg_csr_3453 = _RAND_3453[31:0];
  _RAND_3454 = {1{`RANDOM}};
  reg_csr_3454 = _RAND_3454[31:0];
  _RAND_3455 = {1{`RANDOM}};
  reg_csr_3455 = _RAND_3455[31:0];
  _RAND_3456 = {1{`RANDOM}};
  reg_csr_3456 = _RAND_3456[31:0];
  _RAND_3457 = {1{`RANDOM}};
  reg_csr_3457 = _RAND_3457[31:0];
  _RAND_3458 = {1{`RANDOM}};
  reg_csr_3458 = _RAND_3458[31:0];
  _RAND_3459 = {1{`RANDOM}};
  reg_csr_3459 = _RAND_3459[31:0];
  _RAND_3460 = {1{`RANDOM}};
  reg_csr_3460 = _RAND_3460[31:0];
  _RAND_3461 = {1{`RANDOM}};
  reg_csr_3461 = _RAND_3461[31:0];
  _RAND_3462 = {1{`RANDOM}};
  reg_csr_3462 = _RAND_3462[31:0];
  _RAND_3463 = {1{`RANDOM}};
  reg_csr_3463 = _RAND_3463[31:0];
  _RAND_3464 = {1{`RANDOM}};
  reg_csr_3464 = _RAND_3464[31:0];
  _RAND_3465 = {1{`RANDOM}};
  reg_csr_3465 = _RAND_3465[31:0];
  _RAND_3466 = {1{`RANDOM}};
  reg_csr_3466 = _RAND_3466[31:0];
  _RAND_3467 = {1{`RANDOM}};
  reg_csr_3467 = _RAND_3467[31:0];
  _RAND_3468 = {1{`RANDOM}};
  reg_csr_3468 = _RAND_3468[31:0];
  _RAND_3469 = {1{`RANDOM}};
  reg_csr_3469 = _RAND_3469[31:0];
  _RAND_3470 = {1{`RANDOM}};
  reg_csr_3470 = _RAND_3470[31:0];
  _RAND_3471 = {1{`RANDOM}};
  reg_csr_3471 = _RAND_3471[31:0];
  _RAND_3472 = {1{`RANDOM}};
  reg_csr_3472 = _RAND_3472[31:0];
  _RAND_3473 = {1{`RANDOM}};
  reg_csr_3473 = _RAND_3473[31:0];
  _RAND_3474 = {1{`RANDOM}};
  reg_csr_3474 = _RAND_3474[31:0];
  _RAND_3475 = {1{`RANDOM}};
  reg_csr_3475 = _RAND_3475[31:0];
  _RAND_3476 = {1{`RANDOM}};
  reg_csr_3476 = _RAND_3476[31:0];
  _RAND_3477 = {1{`RANDOM}};
  reg_csr_3477 = _RAND_3477[31:0];
  _RAND_3478 = {1{`RANDOM}};
  reg_csr_3478 = _RAND_3478[31:0];
  _RAND_3479 = {1{`RANDOM}};
  reg_csr_3479 = _RAND_3479[31:0];
  _RAND_3480 = {1{`RANDOM}};
  reg_csr_3480 = _RAND_3480[31:0];
  _RAND_3481 = {1{`RANDOM}};
  reg_csr_3481 = _RAND_3481[31:0];
  _RAND_3482 = {1{`RANDOM}};
  reg_csr_3482 = _RAND_3482[31:0];
  _RAND_3483 = {1{`RANDOM}};
  reg_csr_3483 = _RAND_3483[31:0];
  _RAND_3484 = {1{`RANDOM}};
  reg_csr_3484 = _RAND_3484[31:0];
  _RAND_3485 = {1{`RANDOM}};
  reg_csr_3485 = _RAND_3485[31:0];
  _RAND_3486 = {1{`RANDOM}};
  reg_csr_3486 = _RAND_3486[31:0];
  _RAND_3487 = {1{`RANDOM}};
  reg_csr_3487 = _RAND_3487[31:0];
  _RAND_3488 = {1{`RANDOM}};
  reg_csr_3488 = _RAND_3488[31:0];
  _RAND_3489 = {1{`RANDOM}};
  reg_csr_3489 = _RAND_3489[31:0];
  _RAND_3490 = {1{`RANDOM}};
  reg_csr_3490 = _RAND_3490[31:0];
  _RAND_3491 = {1{`RANDOM}};
  reg_csr_3491 = _RAND_3491[31:0];
  _RAND_3492 = {1{`RANDOM}};
  reg_csr_3492 = _RAND_3492[31:0];
  _RAND_3493 = {1{`RANDOM}};
  reg_csr_3493 = _RAND_3493[31:0];
  _RAND_3494 = {1{`RANDOM}};
  reg_csr_3494 = _RAND_3494[31:0];
  _RAND_3495 = {1{`RANDOM}};
  reg_csr_3495 = _RAND_3495[31:0];
  _RAND_3496 = {1{`RANDOM}};
  reg_csr_3496 = _RAND_3496[31:0];
  _RAND_3497 = {1{`RANDOM}};
  reg_csr_3497 = _RAND_3497[31:0];
  _RAND_3498 = {1{`RANDOM}};
  reg_csr_3498 = _RAND_3498[31:0];
  _RAND_3499 = {1{`RANDOM}};
  reg_csr_3499 = _RAND_3499[31:0];
  _RAND_3500 = {1{`RANDOM}};
  reg_csr_3500 = _RAND_3500[31:0];
  _RAND_3501 = {1{`RANDOM}};
  reg_csr_3501 = _RAND_3501[31:0];
  _RAND_3502 = {1{`RANDOM}};
  reg_csr_3502 = _RAND_3502[31:0];
  _RAND_3503 = {1{`RANDOM}};
  reg_csr_3503 = _RAND_3503[31:0];
  _RAND_3504 = {1{`RANDOM}};
  reg_csr_3504 = _RAND_3504[31:0];
  _RAND_3505 = {1{`RANDOM}};
  reg_csr_3505 = _RAND_3505[31:0];
  _RAND_3506 = {1{`RANDOM}};
  reg_csr_3506 = _RAND_3506[31:0];
  _RAND_3507 = {1{`RANDOM}};
  reg_csr_3507 = _RAND_3507[31:0];
  _RAND_3508 = {1{`RANDOM}};
  reg_csr_3508 = _RAND_3508[31:0];
  _RAND_3509 = {1{`RANDOM}};
  reg_csr_3509 = _RAND_3509[31:0];
  _RAND_3510 = {1{`RANDOM}};
  reg_csr_3510 = _RAND_3510[31:0];
  _RAND_3511 = {1{`RANDOM}};
  reg_csr_3511 = _RAND_3511[31:0];
  _RAND_3512 = {1{`RANDOM}};
  reg_csr_3512 = _RAND_3512[31:0];
  _RAND_3513 = {1{`RANDOM}};
  reg_csr_3513 = _RAND_3513[31:0];
  _RAND_3514 = {1{`RANDOM}};
  reg_csr_3514 = _RAND_3514[31:0];
  _RAND_3515 = {1{`RANDOM}};
  reg_csr_3515 = _RAND_3515[31:0];
  _RAND_3516 = {1{`RANDOM}};
  reg_csr_3516 = _RAND_3516[31:0];
  _RAND_3517 = {1{`RANDOM}};
  reg_csr_3517 = _RAND_3517[31:0];
  _RAND_3518 = {1{`RANDOM}};
  reg_csr_3518 = _RAND_3518[31:0];
  _RAND_3519 = {1{`RANDOM}};
  reg_csr_3519 = _RAND_3519[31:0];
  _RAND_3520 = {1{`RANDOM}};
  reg_csr_3520 = _RAND_3520[31:0];
  _RAND_3521 = {1{`RANDOM}};
  reg_csr_3521 = _RAND_3521[31:0];
  _RAND_3522 = {1{`RANDOM}};
  reg_csr_3522 = _RAND_3522[31:0];
  _RAND_3523 = {1{`RANDOM}};
  reg_csr_3523 = _RAND_3523[31:0];
  _RAND_3524 = {1{`RANDOM}};
  reg_csr_3524 = _RAND_3524[31:0];
  _RAND_3525 = {1{`RANDOM}};
  reg_csr_3525 = _RAND_3525[31:0];
  _RAND_3526 = {1{`RANDOM}};
  reg_csr_3526 = _RAND_3526[31:0];
  _RAND_3527 = {1{`RANDOM}};
  reg_csr_3527 = _RAND_3527[31:0];
  _RAND_3528 = {1{`RANDOM}};
  reg_csr_3528 = _RAND_3528[31:0];
  _RAND_3529 = {1{`RANDOM}};
  reg_csr_3529 = _RAND_3529[31:0];
  _RAND_3530 = {1{`RANDOM}};
  reg_csr_3530 = _RAND_3530[31:0];
  _RAND_3531 = {1{`RANDOM}};
  reg_csr_3531 = _RAND_3531[31:0];
  _RAND_3532 = {1{`RANDOM}};
  reg_csr_3532 = _RAND_3532[31:0];
  _RAND_3533 = {1{`RANDOM}};
  reg_csr_3533 = _RAND_3533[31:0];
  _RAND_3534 = {1{`RANDOM}};
  reg_csr_3534 = _RAND_3534[31:0];
  _RAND_3535 = {1{`RANDOM}};
  reg_csr_3535 = _RAND_3535[31:0];
  _RAND_3536 = {1{`RANDOM}};
  reg_csr_3536 = _RAND_3536[31:0];
  _RAND_3537 = {1{`RANDOM}};
  reg_csr_3537 = _RAND_3537[31:0];
  _RAND_3538 = {1{`RANDOM}};
  reg_csr_3538 = _RAND_3538[31:0];
  _RAND_3539 = {1{`RANDOM}};
  reg_csr_3539 = _RAND_3539[31:0];
  _RAND_3540 = {1{`RANDOM}};
  reg_csr_3540 = _RAND_3540[31:0];
  _RAND_3541 = {1{`RANDOM}};
  reg_csr_3541 = _RAND_3541[31:0];
  _RAND_3542 = {1{`RANDOM}};
  reg_csr_3542 = _RAND_3542[31:0];
  _RAND_3543 = {1{`RANDOM}};
  reg_csr_3543 = _RAND_3543[31:0];
  _RAND_3544 = {1{`RANDOM}};
  reg_csr_3544 = _RAND_3544[31:0];
  _RAND_3545 = {1{`RANDOM}};
  reg_csr_3545 = _RAND_3545[31:0];
  _RAND_3546 = {1{`RANDOM}};
  reg_csr_3546 = _RAND_3546[31:0];
  _RAND_3547 = {1{`RANDOM}};
  reg_csr_3547 = _RAND_3547[31:0];
  _RAND_3548 = {1{`RANDOM}};
  reg_csr_3548 = _RAND_3548[31:0];
  _RAND_3549 = {1{`RANDOM}};
  reg_csr_3549 = _RAND_3549[31:0];
  _RAND_3550 = {1{`RANDOM}};
  reg_csr_3550 = _RAND_3550[31:0];
  _RAND_3551 = {1{`RANDOM}};
  reg_csr_3551 = _RAND_3551[31:0];
  _RAND_3552 = {1{`RANDOM}};
  reg_csr_3552 = _RAND_3552[31:0];
  _RAND_3553 = {1{`RANDOM}};
  reg_csr_3553 = _RAND_3553[31:0];
  _RAND_3554 = {1{`RANDOM}};
  reg_csr_3554 = _RAND_3554[31:0];
  _RAND_3555 = {1{`RANDOM}};
  reg_csr_3555 = _RAND_3555[31:0];
  _RAND_3556 = {1{`RANDOM}};
  reg_csr_3556 = _RAND_3556[31:0];
  _RAND_3557 = {1{`RANDOM}};
  reg_csr_3557 = _RAND_3557[31:0];
  _RAND_3558 = {1{`RANDOM}};
  reg_csr_3558 = _RAND_3558[31:0];
  _RAND_3559 = {1{`RANDOM}};
  reg_csr_3559 = _RAND_3559[31:0];
  _RAND_3560 = {1{`RANDOM}};
  reg_csr_3560 = _RAND_3560[31:0];
  _RAND_3561 = {1{`RANDOM}};
  reg_csr_3561 = _RAND_3561[31:0];
  _RAND_3562 = {1{`RANDOM}};
  reg_csr_3562 = _RAND_3562[31:0];
  _RAND_3563 = {1{`RANDOM}};
  reg_csr_3563 = _RAND_3563[31:0];
  _RAND_3564 = {1{`RANDOM}};
  reg_csr_3564 = _RAND_3564[31:0];
  _RAND_3565 = {1{`RANDOM}};
  reg_csr_3565 = _RAND_3565[31:0];
  _RAND_3566 = {1{`RANDOM}};
  reg_csr_3566 = _RAND_3566[31:0];
  _RAND_3567 = {1{`RANDOM}};
  reg_csr_3567 = _RAND_3567[31:0];
  _RAND_3568 = {1{`RANDOM}};
  reg_csr_3568 = _RAND_3568[31:0];
  _RAND_3569 = {1{`RANDOM}};
  reg_csr_3569 = _RAND_3569[31:0];
  _RAND_3570 = {1{`RANDOM}};
  reg_csr_3570 = _RAND_3570[31:0];
  _RAND_3571 = {1{`RANDOM}};
  reg_csr_3571 = _RAND_3571[31:0];
  _RAND_3572 = {1{`RANDOM}};
  reg_csr_3572 = _RAND_3572[31:0];
  _RAND_3573 = {1{`RANDOM}};
  reg_csr_3573 = _RAND_3573[31:0];
  _RAND_3574 = {1{`RANDOM}};
  reg_csr_3574 = _RAND_3574[31:0];
  _RAND_3575 = {1{`RANDOM}};
  reg_csr_3575 = _RAND_3575[31:0];
  _RAND_3576 = {1{`RANDOM}};
  reg_csr_3576 = _RAND_3576[31:0];
  _RAND_3577 = {1{`RANDOM}};
  reg_csr_3577 = _RAND_3577[31:0];
  _RAND_3578 = {1{`RANDOM}};
  reg_csr_3578 = _RAND_3578[31:0];
  _RAND_3579 = {1{`RANDOM}};
  reg_csr_3579 = _RAND_3579[31:0];
  _RAND_3580 = {1{`RANDOM}};
  reg_csr_3580 = _RAND_3580[31:0];
  _RAND_3581 = {1{`RANDOM}};
  reg_csr_3581 = _RAND_3581[31:0];
  _RAND_3582 = {1{`RANDOM}};
  reg_csr_3582 = _RAND_3582[31:0];
  _RAND_3583 = {1{`RANDOM}};
  reg_csr_3583 = _RAND_3583[31:0];
  _RAND_3584 = {1{`RANDOM}};
  reg_csr_3584 = _RAND_3584[31:0];
  _RAND_3585 = {1{`RANDOM}};
  reg_csr_3585 = _RAND_3585[31:0];
  _RAND_3586 = {1{`RANDOM}};
  reg_csr_3586 = _RAND_3586[31:0];
  _RAND_3587 = {1{`RANDOM}};
  reg_csr_3587 = _RAND_3587[31:0];
  _RAND_3588 = {1{`RANDOM}};
  reg_csr_3588 = _RAND_3588[31:0];
  _RAND_3589 = {1{`RANDOM}};
  reg_csr_3589 = _RAND_3589[31:0];
  _RAND_3590 = {1{`RANDOM}};
  reg_csr_3590 = _RAND_3590[31:0];
  _RAND_3591 = {1{`RANDOM}};
  reg_csr_3591 = _RAND_3591[31:0];
  _RAND_3592 = {1{`RANDOM}};
  reg_csr_3592 = _RAND_3592[31:0];
  _RAND_3593 = {1{`RANDOM}};
  reg_csr_3593 = _RAND_3593[31:0];
  _RAND_3594 = {1{`RANDOM}};
  reg_csr_3594 = _RAND_3594[31:0];
  _RAND_3595 = {1{`RANDOM}};
  reg_csr_3595 = _RAND_3595[31:0];
  _RAND_3596 = {1{`RANDOM}};
  reg_csr_3596 = _RAND_3596[31:0];
  _RAND_3597 = {1{`RANDOM}};
  reg_csr_3597 = _RAND_3597[31:0];
  _RAND_3598 = {1{`RANDOM}};
  reg_csr_3598 = _RAND_3598[31:0];
  _RAND_3599 = {1{`RANDOM}};
  reg_csr_3599 = _RAND_3599[31:0];
  _RAND_3600 = {1{`RANDOM}};
  reg_csr_3600 = _RAND_3600[31:0];
  _RAND_3601 = {1{`RANDOM}};
  reg_csr_3601 = _RAND_3601[31:0];
  _RAND_3602 = {1{`RANDOM}};
  reg_csr_3602 = _RAND_3602[31:0];
  _RAND_3603 = {1{`RANDOM}};
  reg_csr_3603 = _RAND_3603[31:0];
  _RAND_3604 = {1{`RANDOM}};
  reg_csr_3604 = _RAND_3604[31:0];
  _RAND_3605 = {1{`RANDOM}};
  reg_csr_3605 = _RAND_3605[31:0];
  _RAND_3606 = {1{`RANDOM}};
  reg_csr_3606 = _RAND_3606[31:0];
  _RAND_3607 = {1{`RANDOM}};
  reg_csr_3607 = _RAND_3607[31:0];
  _RAND_3608 = {1{`RANDOM}};
  reg_csr_3608 = _RAND_3608[31:0];
  _RAND_3609 = {1{`RANDOM}};
  reg_csr_3609 = _RAND_3609[31:0];
  _RAND_3610 = {1{`RANDOM}};
  reg_csr_3610 = _RAND_3610[31:0];
  _RAND_3611 = {1{`RANDOM}};
  reg_csr_3611 = _RAND_3611[31:0];
  _RAND_3612 = {1{`RANDOM}};
  reg_csr_3612 = _RAND_3612[31:0];
  _RAND_3613 = {1{`RANDOM}};
  reg_csr_3613 = _RAND_3613[31:0];
  _RAND_3614 = {1{`RANDOM}};
  reg_csr_3614 = _RAND_3614[31:0];
  _RAND_3615 = {1{`RANDOM}};
  reg_csr_3615 = _RAND_3615[31:0];
  _RAND_3616 = {1{`RANDOM}};
  reg_csr_3616 = _RAND_3616[31:0];
  _RAND_3617 = {1{`RANDOM}};
  reg_csr_3617 = _RAND_3617[31:0];
  _RAND_3618 = {1{`RANDOM}};
  reg_csr_3618 = _RAND_3618[31:0];
  _RAND_3619 = {1{`RANDOM}};
  reg_csr_3619 = _RAND_3619[31:0];
  _RAND_3620 = {1{`RANDOM}};
  reg_csr_3620 = _RAND_3620[31:0];
  _RAND_3621 = {1{`RANDOM}};
  reg_csr_3621 = _RAND_3621[31:0];
  _RAND_3622 = {1{`RANDOM}};
  reg_csr_3622 = _RAND_3622[31:0];
  _RAND_3623 = {1{`RANDOM}};
  reg_csr_3623 = _RAND_3623[31:0];
  _RAND_3624 = {1{`RANDOM}};
  reg_csr_3624 = _RAND_3624[31:0];
  _RAND_3625 = {1{`RANDOM}};
  reg_csr_3625 = _RAND_3625[31:0];
  _RAND_3626 = {1{`RANDOM}};
  reg_csr_3626 = _RAND_3626[31:0];
  _RAND_3627 = {1{`RANDOM}};
  reg_csr_3627 = _RAND_3627[31:0];
  _RAND_3628 = {1{`RANDOM}};
  reg_csr_3628 = _RAND_3628[31:0];
  _RAND_3629 = {1{`RANDOM}};
  reg_csr_3629 = _RAND_3629[31:0];
  _RAND_3630 = {1{`RANDOM}};
  reg_csr_3630 = _RAND_3630[31:0];
  _RAND_3631 = {1{`RANDOM}};
  reg_csr_3631 = _RAND_3631[31:0];
  _RAND_3632 = {1{`RANDOM}};
  reg_csr_3632 = _RAND_3632[31:0];
  _RAND_3633 = {1{`RANDOM}};
  reg_csr_3633 = _RAND_3633[31:0];
  _RAND_3634 = {1{`RANDOM}};
  reg_csr_3634 = _RAND_3634[31:0];
  _RAND_3635 = {1{`RANDOM}};
  reg_csr_3635 = _RAND_3635[31:0];
  _RAND_3636 = {1{`RANDOM}};
  reg_csr_3636 = _RAND_3636[31:0];
  _RAND_3637 = {1{`RANDOM}};
  reg_csr_3637 = _RAND_3637[31:0];
  _RAND_3638 = {1{`RANDOM}};
  reg_csr_3638 = _RAND_3638[31:0];
  _RAND_3639 = {1{`RANDOM}};
  reg_csr_3639 = _RAND_3639[31:0];
  _RAND_3640 = {1{`RANDOM}};
  reg_csr_3640 = _RAND_3640[31:0];
  _RAND_3641 = {1{`RANDOM}};
  reg_csr_3641 = _RAND_3641[31:0];
  _RAND_3642 = {1{`RANDOM}};
  reg_csr_3642 = _RAND_3642[31:0];
  _RAND_3643 = {1{`RANDOM}};
  reg_csr_3643 = _RAND_3643[31:0];
  _RAND_3644 = {1{`RANDOM}};
  reg_csr_3644 = _RAND_3644[31:0];
  _RAND_3645 = {1{`RANDOM}};
  reg_csr_3645 = _RAND_3645[31:0];
  _RAND_3646 = {1{`RANDOM}};
  reg_csr_3646 = _RAND_3646[31:0];
  _RAND_3647 = {1{`RANDOM}};
  reg_csr_3647 = _RAND_3647[31:0];
  _RAND_3648 = {1{`RANDOM}};
  reg_csr_3648 = _RAND_3648[31:0];
  _RAND_3649 = {1{`RANDOM}};
  reg_csr_3649 = _RAND_3649[31:0];
  _RAND_3650 = {1{`RANDOM}};
  reg_csr_3650 = _RAND_3650[31:0];
  _RAND_3651 = {1{`RANDOM}};
  reg_csr_3651 = _RAND_3651[31:0];
  _RAND_3652 = {1{`RANDOM}};
  reg_csr_3652 = _RAND_3652[31:0];
  _RAND_3653 = {1{`RANDOM}};
  reg_csr_3653 = _RAND_3653[31:0];
  _RAND_3654 = {1{`RANDOM}};
  reg_csr_3654 = _RAND_3654[31:0];
  _RAND_3655 = {1{`RANDOM}};
  reg_csr_3655 = _RAND_3655[31:0];
  _RAND_3656 = {1{`RANDOM}};
  reg_csr_3656 = _RAND_3656[31:0];
  _RAND_3657 = {1{`RANDOM}};
  reg_csr_3657 = _RAND_3657[31:0];
  _RAND_3658 = {1{`RANDOM}};
  reg_csr_3658 = _RAND_3658[31:0];
  _RAND_3659 = {1{`RANDOM}};
  reg_csr_3659 = _RAND_3659[31:0];
  _RAND_3660 = {1{`RANDOM}};
  reg_csr_3660 = _RAND_3660[31:0];
  _RAND_3661 = {1{`RANDOM}};
  reg_csr_3661 = _RAND_3661[31:0];
  _RAND_3662 = {1{`RANDOM}};
  reg_csr_3662 = _RAND_3662[31:0];
  _RAND_3663 = {1{`RANDOM}};
  reg_csr_3663 = _RAND_3663[31:0];
  _RAND_3664 = {1{`RANDOM}};
  reg_csr_3664 = _RAND_3664[31:0];
  _RAND_3665 = {1{`RANDOM}};
  reg_csr_3665 = _RAND_3665[31:0];
  _RAND_3666 = {1{`RANDOM}};
  reg_csr_3666 = _RAND_3666[31:0];
  _RAND_3667 = {1{`RANDOM}};
  reg_csr_3667 = _RAND_3667[31:0];
  _RAND_3668 = {1{`RANDOM}};
  reg_csr_3668 = _RAND_3668[31:0];
  _RAND_3669 = {1{`RANDOM}};
  reg_csr_3669 = _RAND_3669[31:0];
  _RAND_3670 = {1{`RANDOM}};
  reg_csr_3670 = _RAND_3670[31:0];
  _RAND_3671 = {1{`RANDOM}};
  reg_csr_3671 = _RAND_3671[31:0];
  _RAND_3672 = {1{`RANDOM}};
  reg_csr_3672 = _RAND_3672[31:0];
  _RAND_3673 = {1{`RANDOM}};
  reg_csr_3673 = _RAND_3673[31:0];
  _RAND_3674 = {1{`RANDOM}};
  reg_csr_3674 = _RAND_3674[31:0];
  _RAND_3675 = {1{`RANDOM}};
  reg_csr_3675 = _RAND_3675[31:0];
  _RAND_3676 = {1{`RANDOM}};
  reg_csr_3676 = _RAND_3676[31:0];
  _RAND_3677 = {1{`RANDOM}};
  reg_csr_3677 = _RAND_3677[31:0];
  _RAND_3678 = {1{`RANDOM}};
  reg_csr_3678 = _RAND_3678[31:0];
  _RAND_3679 = {1{`RANDOM}};
  reg_csr_3679 = _RAND_3679[31:0];
  _RAND_3680 = {1{`RANDOM}};
  reg_csr_3680 = _RAND_3680[31:0];
  _RAND_3681 = {1{`RANDOM}};
  reg_csr_3681 = _RAND_3681[31:0];
  _RAND_3682 = {1{`RANDOM}};
  reg_csr_3682 = _RAND_3682[31:0];
  _RAND_3683 = {1{`RANDOM}};
  reg_csr_3683 = _RAND_3683[31:0];
  _RAND_3684 = {1{`RANDOM}};
  reg_csr_3684 = _RAND_3684[31:0];
  _RAND_3685 = {1{`RANDOM}};
  reg_csr_3685 = _RAND_3685[31:0];
  _RAND_3686 = {1{`RANDOM}};
  reg_csr_3686 = _RAND_3686[31:0];
  _RAND_3687 = {1{`RANDOM}};
  reg_csr_3687 = _RAND_3687[31:0];
  _RAND_3688 = {1{`RANDOM}};
  reg_csr_3688 = _RAND_3688[31:0];
  _RAND_3689 = {1{`RANDOM}};
  reg_csr_3689 = _RAND_3689[31:0];
  _RAND_3690 = {1{`RANDOM}};
  reg_csr_3690 = _RAND_3690[31:0];
  _RAND_3691 = {1{`RANDOM}};
  reg_csr_3691 = _RAND_3691[31:0];
  _RAND_3692 = {1{`RANDOM}};
  reg_csr_3692 = _RAND_3692[31:0];
  _RAND_3693 = {1{`RANDOM}};
  reg_csr_3693 = _RAND_3693[31:0];
  _RAND_3694 = {1{`RANDOM}};
  reg_csr_3694 = _RAND_3694[31:0];
  _RAND_3695 = {1{`RANDOM}};
  reg_csr_3695 = _RAND_3695[31:0];
  _RAND_3696 = {1{`RANDOM}};
  reg_csr_3696 = _RAND_3696[31:0];
  _RAND_3697 = {1{`RANDOM}};
  reg_csr_3697 = _RAND_3697[31:0];
  _RAND_3698 = {1{`RANDOM}};
  reg_csr_3698 = _RAND_3698[31:0];
  _RAND_3699 = {1{`RANDOM}};
  reg_csr_3699 = _RAND_3699[31:0];
  _RAND_3700 = {1{`RANDOM}};
  reg_csr_3700 = _RAND_3700[31:0];
  _RAND_3701 = {1{`RANDOM}};
  reg_csr_3701 = _RAND_3701[31:0];
  _RAND_3702 = {1{`RANDOM}};
  reg_csr_3702 = _RAND_3702[31:0];
  _RAND_3703 = {1{`RANDOM}};
  reg_csr_3703 = _RAND_3703[31:0];
  _RAND_3704 = {1{`RANDOM}};
  reg_csr_3704 = _RAND_3704[31:0];
  _RAND_3705 = {1{`RANDOM}};
  reg_csr_3705 = _RAND_3705[31:0];
  _RAND_3706 = {1{`RANDOM}};
  reg_csr_3706 = _RAND_3706[31:0];
  _RAND_3707 = {1{`RANDOM}};
  reg_csr_3707 = _RAND_3707[31:0];
  _RAND_3708 = {1{`RANDOM}};
  reg_csr_3708 = _RAND_3708[31:0];
  _RAND_3709 = {1{`RANDOM}};
  reg_csr_3709 = _RAND_3709[31:0];
  _RAND_3710 = {1{`RANDOM}};
  reg_csr_3710 = _RAND_3710[31:0];
  _RAND_3711 = {1{`RANDOM}};
  reg_csr_3711 = _RAND_3711[31:0];
  _RAND_3712 = {1{`RANDOM}};
  reg_csr_3712 = _RAND_3712[31:0];
  _RAND_3713 = {1{`RANDOM}};
  reg_csr_3713 = _RAND_3713[31:0];
  _RAND_3714 = {1{`RANDOM}};
  reg_csr_3714 = _RAND_3714[31:0];
  _RAND_3715 = {1{`RANDOM}};
  reg_csr_3715 = _RAND_3715[31:0];
  _RAND_3716 = {1{`RANDOM}};
  reg_csr_3716 = _RAND_3716[31:0];
  _RAND_3717 = {1{`RANDOM}};
  reg_csr_3717 = _RAND_3717[31:0];
  _RAND_3718 = {1{`RANDOM}};
  reg_csr_3718 = _RAND_3718[31:0];
  _RAND_3719 = {1{`RANDOM}};
  reg_csr_3719 = _RAND_3719[31:0];
  _RAND_3720 = {1{`RANDOM}};
  reg_csr_3720 = _RAND_3720[31:0];
  _RAND_3721 = {1{`RANDOM}};
  reg_csr_3721 = _RAND_3721[31:0];
  _RAND_3722 = {1{`RANDOM}};
  reg_csr_3722 = _RAND_3722[31:0];
  _RAND_3723 = {1{`RANDOM}};
  reg_csr_3723 = _RAND_3723[31:0];
  _RAND_3724 = {1{`RANDOM}};
  reg_csr_3724 = _RAND_3724[31:0];
  _RAND_3725 = {1{`RANDOM}};
  reg_csr_3725 = _RAND_3725[31:0];
  _RAND_3726 = {1{`RANDOM}};
  reg_csr_3726 = _RAND_3726[31:0];
  _RAND_3727 = {1{`RANDOM}};
  reg_csr_3727 = _RAND_3727[31:0];
  _RAND_3728 = {1{`RANDOM}};
  reg_csr_3728 = _RAND_3728[31:0];
  _RAND_3729 = {1{`RANDOM}};
  reg_csr_3729 = _RAND_3729[31:0];
  _RAND_3730 = {1{`RANDOM}};
  reg_csr_3730 = _RAND_3730[31:0];
  _RAND_3731 = {1{`RANDOM}};
  reg_csr_3731 = _RAND_3731[31:0];
  _RAND_3732 = {1{`RANDOM}};
  reg_csr_3732 = _RAND_3732[31:0];
  _RAND_3733 = {1{`RANDOM}};
  reg_csr_3733 = _RAND_3733[31:0];
  _RAND_3734 = {1{`RANDOM}};
  reg_csr_3734 = _RAND_3734[31:0];
  _RAND_3735 = {1{`RANDOM}};
  reg_csr_3735 = _RAND_3735[31:0];
  _RAND_3736 = {1{`RANDOM}};
  reg_csr_3736 = _RAND_3736[31:0];
  _RAND_3737 = {1{`RANDOM}};
  reg_csr_3737 = _RAND_3737[31:0];
  _RAND_3738 = {1{`RANDOM}};
  reg_csr_3738 = _RAND_3738[31:0];
  _RAND_3739 = {1{`RANDOM}};
  reg_csr_3739 = _RAND_3739[31:0];
  _RAND_3740 = {1{`RANDOM}};
  reg_csr_3740 = _RAND_3740[31:0];
  _RAND_3741 = {1{`RANDOM}};
  reg_csr_3741 = _RAND_3741[31:0];
  _RAND_3742 = {1{`RANDOM}};
  reg_csr_3742 = _RAND_3742[31:0];
  _RAND_3743 = {1{`RANDOM}};
  reg_csr_3743 = _RAND_3743[31:0];
  _RAND_3744 = {1{`RANDOM}};
  reg_csr_3744 = _RAND_3744[31:0];
  _RAND_3745 = {1{`RANDOM}};
  reg_csr_3745 = _RAND_3745[31:0];
  _RAND_3746 = {1{`RANDOM}};
  reg_csr_3746 = _RAND_3746[31:0];
  _RAND_3747 = {1{`RANDOM}};
  reg_csr_3747 = _RAND_3747[31:0];
  _RAND_3748 = {1{`RANDOM}};
  reg_csr_3748 = _RAND_3748[31:0];
  _RAND_3749 = {1{`RANDOM}};
  reg_csr_3749 = _RAND_3749[31:0];
  _RAND_3750 = {1{`RANDOM}};
  reg_csr_3750 = _RAND_3750[31:0];
  _RAND_3751 = {1{`RANDOM}};
  reg_csr_3751 = _RAND_3751[31:0];
  _RAND_3752 = {1{`RANDOM}};
  reg_csr_3752 = _RAND_3752[31:0];
  _RAND_3753 = {1{`RANDOM}};
  reg_csr_3753 = _RAND_3753[31:0];
  _RAND_3754 = {1{`RANDOM}};
  reg_csr_3754 = _RAND_3754[31:0];
  _RAND_3755 = {1{`RANDOM}};
  reg_csr_3755 = _RAND_3755[31:0];
  _RAND_3756 = {1{`RANDOM}};
  reg_csr_3756 = _RAND_3756[31:0];
  _RAND_3757 = {1{`RANDOM}};
  reg_csr_3757 = _RAND_3757[31:0];
  _RAND_3758 = {1{`RANDOM}};
  reg_csr_3758 = _RAND_3758[31:0];
  _RAND_3759 = {1{`RANDOM}};
  reg_csr_3759 = _RAND_3759[31:0];
  _RAND_3760 = {1{`RANDOM}};
  reg_csr_3760 = _RAND_3760[31:0];
  _RAND_3761 = {1{`RANDOM}};
  reg_csr_3761 = _RAND_3761[31:0];
  _RAND_3762 = {1{`RANDOM}};
  reg_csr_3762 = _RAND_3762[31:0];
  _RAND_3763 = {1{`RANDOM}};
  reg_csr_3763 = _RAND_3763[31:0];
  _RAND_3764 = {1{`RANDOM}};
  reg_csr_3764 = _RAND_3764[31:0];
  _RAND_3765 = {1{`RANDOM}};
  reg_csr_3765 = _RAND_3765[31:0];
  _RAND_3766 = {1{`RANDOM}};
  reg_csr_3766 = _RAND_3766[31:0];
  _RAND_3767 = {1{`RANDOM}};
  reg_csr_3767 = _RAND_3767[31:0];
  _RAND_3768 = {1{`RANDOM}};
  reg_csr_3768 = _RAND_3768[31:0];
  _RAND_3769 = {1{`RANDOM}};
  reg_csr_3769 = _RAND_3769[31:0];
  _RAND_3770 = {1{`RANDOM}};
  reg_csr_3770 = _RAND_3770[31:0];
  _RAND_3771 = {1{`RANDOM}};
  reg_csr_3771 = _RAND_3771[31:0];
  _RAND_3772 = {1{`RANDOM}};
  reg_csr_3772 = _RAND_3772[31:0];
  _RAND_3773 = {1{`RANDOM}};
  reg_csr_3773 = _RAND_3773[31:0];
  _RAND_3774 = {1{`RANDOM}};
  reg_csr_3774 = _RAND_3774[31:0];
  _RAND_3775 = {1{`RANDOM}};
  reg_csr_3775 = _RAND_3775[31:0];
  _RAND_3776 = {1{`RANDOM}};
  reg_csr_3776 = _RAND_3776[31:0];
  _RAND_3777 = {1{`RANDOM}};
  reg_csr_3777 = _RAND_3777[31:0];
  _RAND_3778 = {1{`RANDOM}};
  reg_csr_3778 = _RAND_3778[31:0];
  _RAND_3779 = {1{`RANDOM}};
  reg_csr_3779 = _RAND_3779[31:0];
  _RAND_3780 = {1{`RANDOM}};
  reg_csr_3780 = _RAND_3780[31:0];
  _RAND_3781 = {1{`RANDOM}};
  reg_csr_3781 = _RAND_3781[31:0];
  _RAND_3782 = {1{`RANDOM}};
  reg_csr_3782 = _RAND_3782[31:0];
  _RAND_3783 = {1{`RANDOM}};
  reg_csr_3783 = _RAND_3783[31:0];
  _RAND_3784 = {1{`RANDOM}};
  reg_csr_3784 = _RAND_3784[31:0];
  _RAND_3785 = {1{`RANDOM}};
  reg_csr_3785 = _RAND_3785[31:0];
  _RAND_3786 = {1{`RANDOM}};
  reg_csr_3786 = _RAND_3786[31:0];
  _RAND_3787 = {1{`RANDOM}};
  reg_csr_3787 = _RAND_3787[31:0];
  _RAND_3788 = {1{`RANDOM}};
  reg_csr_3788 = _RAND_3788[31:0];
  _RAND_3789 = {1{`RANDOM}};
  reg_csr_3789 = _RAND_3789[31:0];
  _RAND_3790 = {1{`RANDOM}};
  reg_csr_3790 = _RAND_3790[31:0];
  _RAND_3791 = {1{`RANDOM}};
  reg_csr_3791 = _RAND_3791[31:0];
  _RAND_3792 = {1{`RANDOM}};
  reg_csr_3792 = _RAND_3792[31:0];
  _RAND_3793 = {1{`RANDOM}};
  reg_csr_3793 = _RAND_3793[31:0];
  _RAND_3794 = {1{`RANDOM}};
  reg_csr_3794 = _RAND_3794[31:0];
  _RAND_3795 = {1{`RANDOM}};
  reg_csr_3795 = _RAND_3795[31:0];
  _RAND_3796 = {1{`RANDOM}};
  reg_csr_3796 = _RAND_3796[31:0];
  _RAND_3797 = {1{`RANDOM}};
  reg_csr_3797 = _RAND_3797[31:0];
  _RAND_3798 = {1{`RANDOM}};
  reg_csr_3798 = _RAND_3798[31:0];
  _RAND_3799 = {1{`RANDOM}};
  reg_csr_3799 = _RAND_3799[31:0];
  _RAND_3800 = {1{`RANDOM}};
  reg_csr_3800 = _RAND_3800[31:0];
  _RAND_3801 = {1{`RANDOM}};
  reg_csr_3801 = _RAND_3801[31:0];
  _RAND_3802 = {1{`RANDOM}};
  reg_csr_3802 = _RAND_3802[31:0];
  _RAND_3803 = {1{`RANDOM}};
  reg_csr_3803 = _RAND_3803[31:0];
  _RAND_3804 = {1{`RANDOM}};
  reg_csr_3804 = _RAND_3804[31:0];
  _RAND_3805 = {1{`RANDOM}};
  reg_csr_3805 = _RAND_3805[31:0];
  _RAND_3806 = {1{`RANDOM}};
  reg_csr_3806 = _RAND_3806[31:0];
  _RAND_3807 = {1{`RANDOM}};
  reg_csr_3807 = _RAND_3807[31:0];
  _RAND_3808 = {1{`RANDOM}};
  reg_csr_3808 = _RAND_3808[31:0];
  _RAND_3809 = {1{`RANDOM}};
  reg_csr_3809 = _RAND_3809[31:0];
  _RAND_3810 = {1{`RANDOM}};
  reg_csr_3810 = _RAND_3810[31:0];
  _RAND_3811 = {1{`RANDOM}};
  reg_csr_3811 = _RAND_3811[31:0];
  _RAND_3812 = {1{`RANDOM}};
  reg_csr_3812 = _RAND_3812[31:0];
  _RAND_3813 = {1{`RANDOM}};
  reg_csr_3813 = _RAND_3813[31:0];
  _RAND_3814 = {1{`RANDOM}};
  reg_csr_3814 = _RAND_3814[31:0];
  _RAND_3815 = {1{`RANDOM}};
  reg_csr_3815 = _RAND_3815[31:0];
  _RAND_3816 = {1{`RANDOM}};
  reg_csr_3816 = _RAND_3816[31:0];
  _RAND_3817 = {1{`RANDOM}};
  reg_csr_3817 = _RAND_3817[31:0];
  _RAND_3818 = {1{`RANDOM}};
  reg_csr_3818 = _RAND_3818[31:0];
  _RAND_3819 = {1{`RANDOM}};
  reg_csr_3819 = _RAND_3819[31:0];
  _RAND_3820 = {1{`RANDOM}};
  reg_csr_3820 = _RAND_3820[31:0];
  _RAND_3821 = {1{`RANDOM}};
  reg_csr_3821 = _RAND_3821[31:0];
  _RAND_3822 = {1{`RANDOM}};
  reg_csr_3822 = _RAND_3822[31:0];
  _RAND_3823 = {1{`RANDOM}};
  reg_csr_3823 = _RAND_3823[31:0];
  _RAND_3824 = {1{`RANDOM}};
  reg_csr_3824 = _RAND_3824[31:0];
  _RAND_3825 = {1{`RANDOM}};
  reg_csr_3825 = _RAND_3825[31:0];
  _RAND_3826 = {1{`RANDOM}};
  reg_csr_3826 = _RAND_3826[31:0];
  _RAND_3827 = {1{`RANDOM}};
  reg_csr_3827 = _RAND_3827[31:0];
  _RAND_3828 = {1{`RANDOM}};
  reg_csr_3828 = _RAND_3828[31:0];
  _RAND_3829 = {1{`RANDOM}};
  reg_csr_3829 = _RAND_3829[31:0];
  _RAND_3830 = {1{`RANDOM}};
  reg_csr_3830 = _RAND_3830[31:0];
  _RAND_3831 = {1{`RANDOM}};
  reg_csr_3831 = _RAND_3831[31:0];
  _RAND_3832 = {1{`RANDOM}};
  reg_csr_3832 = _RAND_3832[31:0];
  _RAND_3833 = {1{`RANDOM}};
  reg_csr_3833 = _RAND_3833[31:0];
  _RAND_3834 = {1{`RANDOM}};
  reg_csr_3834 = _RAND_3834[31:0];
  _RAND_3835 = {1{`RANDOM}};
  reg_csr_3835 = _RAND_3835[31:0];
  _RAND_3836 = {1{`RANDOM}};
  reg_csr_3836 = _RAND_3836[31:0];
  _RAND_3837 = {1{`RANDOM}};
  reg_csr_3837 = _RAND_3837[31:0];
  _RAND_3838 = {1{`RANDOM}};
  reg_csr_3838 = _RAND_3838[31:0];
  _RAND_3839 = {1{`RANDOM}};
  reg_csr_3839 = _RAND_3839[31:0];
  _RAND_3840 = {1{`RANDOM}};
  reg_csr_3840 = _RAND_3840[31:0];
  _RAND_3841 = {1{`RANDOM}};
  reg_csr_3841 = _RAND_3841[31:0];
  _RAND_3842 = {1{`RANDOM}};
  reg_csr_3842 = _RAND_3842[31:0];
  _RAND_3843 = {1{`RANDOM}};
  reg_csr_3843 = _RAND_3843[31:0];
  _RAND_3844 = {1{`RANDOM}};
  reg_csr_3844 = _RAND_3844[31:0];
  _RAND_3845 = {1{`RANDOM}};
  reg_csr_3845 = _RAND_3845[31:0];
  _RAND_3846 = {1{`RANDOM}};
  reg_csr_3846 = _RAND_3846[31:0];
  _RAND_3847 = {1{`RANDOM}};
  reg_csr_3847 = _RAND_3847[31:0];
  _RAND_3848 = {1{`RANDOM}};
  reg_csr_3848 = _RAND_3848[31:0];
  _RAND_3849 = {1{`RANDOM}};
  reg_csr_3849 = _RAND_3849[31:0];
  _RAND_3850 = {1{`RANDOM}};
  reg_csr_3850 = _RAND_3850[31:0];
  _RAND_3851 = {1{`RANDOM}};
  reg_csr_3851 = _RAND_3851[31:0];
  _RAND_3852 = {1{`RANDOM}};
  reg_csr_3852 = _RAND_3852[31:0];
  _RAND_3853 = {1{`RANDOM}};
  reg_csr_3853 = _RAND_3853[31:0];
  _RAND_3854 = {1{`RANDOM}};
  reg_csr_3854 = _RAND_3854[31:0];
  _RAND_3855 = {1{`RANDOM}};
  reg_csr_3855 = _RAND_3855[31:0];
  _RAND_3856 = {1{`RANDOM}};
  reg_csr_3856 = _RAND_3856[31:0];
  _RAND_3857 = {1{`RANDOM}};
  reg_csr_3857 = _RAND_3857[31:0];
  _RAND_3858 = {1{`RANDOM}};
  reg_csr_3858 = _RAND_3858[31:0];
  _RAND_3859 = {1{`RANDOM}};
  reg_csr_3859 = _RAND_3859[31:0];
  _RAND_3860 = {1{`RANDOM}};
  reg_csr_3860 = _RAND_3860[31:0];
  _RAND_3861 = {1{`RANDOM}};
  reg_csr_3861 = _RAND_3861[31:0];
  _RAND_3862 = {1{`RANDOM}};
  reg_csr_3862 = _RAND_3862[31:0];
  _RAND_3863 = {1{`RANDOM}};
  reg_csr_3863 = _RAND_3863[31:0];
  _RAND_3864 = {1{`RANDOM}};
  reg_csr_3864 = _RAND_3864[31:0];
  _RAND_3865 = {1{`RANDOM}};
  reg_csr_3865 = _RAND_3865[31:0];
  _RAND_3866 = {1{`RANDOM}};
  reg_csr_3866 = _RAND_3866[31:0];
  _RAND_3867 = {1{`RANDOM}};
  reg_csr_3867 = _RAND_3867[31:0];
  _RAND_3868 = {1{`RANDOM}};
  reg_csr_3868 = _RAND_3868[31:0];
  _RAND_3869 = {1{`RANDOM}};
  reg_csr_3869 = _RAND_3869[31:0];
  _RAND_3870 = {1{`RANDOM}};
  reg_csr_3870 = _RAND_3870[31:0];
  _RAND_3871 = {1{`RANDOM}};
  reg_csr_3871 = _RAND_3871[31:0];
  _RAND_3872 = {1{`RANDOM}};
  reg_csr_3872 = _RAND_3872[31:0];
  _RAND_3873 = {1{`RANDOM}};
  reg_csr_3873 = _RAND_3873[31:0];
  _RAND_3874 = {1{`RANDOM}};
  reg_csr_3874 = _RAND_3874[31:0];
  _RAND_3875 = {1{`RANDOM}};
  reg_csr_3875 = _RAND_3875[31:0];
  _RAND_3876 = {1{`RANDOM}};
  reg_csr_3876 = _RAND_3876[31:0];
  _RAND_3877 = {1{`RANDOM}};
  reg_csr_3877 = _RAND_3877[31:0];
  _RAND_3878 = {1{`RANDOM}};
  reg_csr_3878 = _RAND_3878[31:0];
  _RAND_3879 = {1{`RANDOM}};
  reg_csr_3879 = _RAND_3879[31:0];
  _RAND_3880 = {1{`RANDOM}};
  reg_csr_3880 = _RAND_3880[31:0];
  _RAND_3881 = {1{`RANDOM}};
  reg_csr_3881 = _RAND_3881[31:0];
  _RAND_3882 = {1{`RANDOM}};
  reg_csr_3882 = _RAND_3882[31:0];
  _RAND_3883 = {1{`RANDOM}};
  reg_csr_3883 = _RAND_3883[31:0];
  _RAND_3884 = {1{`RANDOM}};
  reg_csr_3884 = _RAND_3884[31:0];
  _RAND_3885 = {1{`RANDOM}};
  reg_csr_3885 = _RAND_3885[31:0];
  _RAND_3886 = {1{`RANDOM}};
  reg_csr_3886 = _RAND_3886[31:0];
  _RAND_3887 = {1{`RANDOM}};
  reg_csr_3887 = _RAND_3887[31:0];
  _RAND_3888 = {1{`RANDOM}};
  reg_csr_3888 = _RAND_3888[31:0];
  _RAND_3889 = {1{`RANDOM}};
  reg_csr_3889 = _RAND_3889[31:0];
  _RAND_3890 = {1{`RANDOM}};
  reg_csr_3890 = _RAND_3890[31:0];
  _RAND_3891 = {1{`RANDOM}};
  reg_csr_3891 = _RAND_3891[31:0];
  _RAND_3892 = {1{`RANDOM}};
  reg_csr_3892 = _RAND_3892[31:0];
  _RAND_3893 = {1{`RANDOM}};
  reg_csr_3893 = _RAND_3893[31:0];
  _RAND_3894 = {1{`RANDOM}};
  reg_csr_3894 = _RAND_3894[31:0];
  _RAND_3895 = {1{`RANDOM}};
  reg_csr_3895 = _RAND_3895[31:0];
  _RAND_3896 = {1{`RANDOM}};
  reg_csr_3896 = _RAND_3896[31:0];
  _RAND_3897 = {1{`RANDOM}};
  reg_csr_3897 = _RAND_3897[31:0];
  _RAND_3898 = {1{`RANDOM}};
  reg_csr_3898 = _RAND_3898[31:0];
  _RAND_3899 = {1{`RANDOM}};
  reg_csr_3899 = _RAND_3899[31:0];
  _RAND_3900 = {1{`RANDOM}};
  reg_csr_3900 = _RAND_3900[31:0];
  _RAND_3901 = {1{`RANDOM}};
  reg_csr_3901 = _RAND_3901[31:0];
  _RAND_3902 = {1{`RANDOM}};
  reg_csr_3902 = _RAND_3902[31:0];
  _RAND_3903 = {1{`RANDOM}};
  reg_csr_3903 = _RAND_3903[31:0];
  _RAND_3904 = {1{`RANDOM}};
  reg_csr_3904 = _RAND_3904[31:0];
  _RAND_3905 = {1{`RANDOM}};
  reg_csr_3905 = _RAND_3905[31:0];
  _RAND_3906 = {1{`RANDOM}};
  reg_csr_3906 = _RAND_3906[31:0];
  _RAND_3907 = {1{`RANDOM}};
  reg_csr_3907 = _RAND_3907[31:0];
  _RAND_3908 = {1{`RANDOM}};
  reg_csr_3908 = _RAND_3908[31:0];
  _RAND_3909 = {1{`RANDOM}};
  reg_csr_3909 = _RAND_3909[31:0];
  _RAND_3910 = {1{`RANDOM}};
  reg_csr_3910 = _RAND_3910[31:0];
  _RAND_3911 = {1{`RANDOM}};
  reg_csr_3911 = _RAND_3911[31:0];
  _RAND_3912 = {1{`RANDOM}};
  reg_csr_3912 = _RAND_3912[31:0];
  _RAND_3913 = {1{`RANDOM}};
  reg_csr_3913 = _RAND_3913[31:0];
  _RAND_3914 = {1{`RANDOM}};
  reg_csr_3914 = _RAND_3914[31:0];
  _RAND_3915 = {1{`RANDOM}};
  reg_csr_3915 = _RAND_3915[31:0];
  _RAND_3916 = {1{`RANDOM}};
  reg_csr_3916 = _RAND_3916[31:0];
  _RAND_3917 = {1{`RANDOM}};
  reg_csr_3917 = _RAND_3917[31:0];
  _RAND_3918 = {1{`RANDOM}};
  reg_csr_3918 = _RAND_3918[31:0];
  _RAND_3919 = {1{`RANDOM}};
  reg_csr_3919 = _RAND_3919[31:0];
  _RAND_3920 = {1{`RANDOM}};
  reg_csr_3920 = _RAND_3920[31:0];
  _RAND_3921 = {1{`RANDOM}};
  reg_csr_3921 = _RAND_3921[31:0];
  _RAND_3922 = {1{`RANDOM}};
  reg_csr_3922 = _RAND_3922[31:0];
  _RAND_3923 = {1{`RANDOM}};
  reg_csr_3923 = _RAND_3923[31:0];
  _RAND_3924 = {1{`RANDOM}};
  reg_csr_3924 = _RAND_3924[31:0];
  _RAND_3925 = {1{`RANDOM}};
  reg_csr_3925 = _RAND_3925[31:0];
  _RAND_3926 = {1{`RANDOM}};
  reg_csr_3926 = _RAND_3926[31:0];
  _RAND_3927 = {1{`RANDOM}};
  reg_csr_3927 = _RAND_3927[31:0];
  _RAND_3928 = {1{`RANDOM}};
  reg_csr_3928 = _RAND_3928[31:0];
  _RAND_3929 = {1{`RANDOM}};
  reg_csr_3929 = _RAND_3929[31:0];
  _RAND_3930 = {1{`RANDOM}};
  reg_csr_3930 = _RAND_3930[31:0];
  _RAND_3931 = {1{`RANDOM}};
  reg_csr_3931 = _RAND_3931[31:0];
  _RAND_3932 = {1{`RANDOM}};
  reg_csr_3932 = _RAND_3932[31:0];
  _RAND_3933 = {1{`RANDOM}};
  reg_csr_3933 = _RAND_3933[31:0];
  _RAND_3934 = {1{`RANDOM}};
  reg_csr_3934 = _RAND_3934[31:0];
  _RAND_3935 = {1{`RANDOM}};
  reg_csr_3935 = _RAND_3935[31:0];
  _RAND_3936 = {1{`RANDOM}};
  reg_csr_3936 = _RAND_3936[31:0];
  _RAND_3937 = {1{`RANDOM}};
  reg_csr_3937 = _RAND_3937[31:0];
  _RAND_3938 = {1{`RANDOM}};
  reg_csr_3938 = _RAND_3938[31:0];
  _RAND_3939 = {1{`RANDOM}};
  reg_csr_3939 = _RAND_3939[31:0];
  _RAND_3940 = {1{`RANDOM}};
  reg_csr_3940 = _RAND_3940[31:0];
  _RAND_3941 = {1{`RANDOM}};
  reg_csr_3941 = _RAND_3941[31:0];
  _RAND_3942 = {1{`RANDOM}};
  reg_csr_3942 = _RAND_3942[31:0];
  _RAND_3943 = {1{`RANDOM}};
  reg_csr_3943 = _RAND_3943[31:0];
  _RAND_3944 = {1{`RANDOM}};
  reg_csr_3944 = _RAND_3944[31:0];
  _RAND_3945 = {1{`RANDOM}};
  reg_csr_3945 = _RAND_3945[31:0];
  _RAND_3946 = {1{`RANDOM}};
  reg_csr_3946 = _RAND_3946[31:0];
  _RAND_3947 = {1{`RANDOM}};
  reg_csr_3947 = _RAND_3947[31:0];
  _RAND_3948 = {1{`RANDOM}};
  reg_csr_3948 = _RAND_3948[31:0];
  _RAND_3949 = {1{`RANDOM}};
  reg_csr_3949 = _RAND_3949[31:0];
  _RAND_3950 = {1{`RANDOM}};
  reg_csr_3950 = _RAND_3950[31:0];
  _RAND_3951 = {1{`RANDOM}};
  reg_csr_3951 = _RAND_3951[31:0];
  _RAND_3952 = {1{`RANDOM}};
  reg_csr_3952 = _RAND_3952[31:0];
  _RAND_3953 = {1{`RANDOM}};
  reg_csr_3953 = _RAND_3953[31:0];
  _RAND_3954 = {1{`RANDOM}};
  reg_csr_3954 = _RAND_3954[31:0];
  _RAND_3955 = {1{`RANDOM}};
  reg_csr_3955 = _RAND_3955[31:0];
  _RAND_3956 = {1{`RANDOM}};
  reg_csr_3956 = _RAND_3956[31:0];
  _RAND_3957 = {1{`RANDOM}};
  reg_csr_3957 = _RAND_3957[31:0];
  _RAND_3958 = {1{`RANDOM}};
  reg_csr_3958 = _RAND_3958[31:0];
  _RAND_3959 = {1{`RANDOM}};
  reg_csr_3959 = _RAND_3959[31:0];
  _RAND_3960 = {1{`RANDOM}};
  reg_csr_3960 = _RAND_3960[31:0];
  _RAND_3961 = {1{`RANDOM}};
  reg_csr_3961 = _RAND_3961[31:0];
  _RAND_3962 = {1{`RANDOM}};
  reg_csr_3962 = _RAND_3962[31:0];
  _RAND_3963 = {1{`RANDOM}};
  reg_csr_3963 = _RAND_3963[31:0];
  _RAND_3964 = {1{`RANDOM}};
  reg_csr_3964 = _RAND_3964[31:0];
  _RAND_3965 = {1{`RANDOM}};
  reg_csr_3965 = _RAND_3965[31:0];
  _RAND_3966 = {1{`RANDOM}};
  reg_csr_3966 = _RAND_3966[31:0];
  _RAND_3967 = {1{`RANDOM}};
  reg_csr_3967 = _RAND_3967[31:0];
  _RAND_3968 = {1{`RANDOM}};
  reg_csr_3968 = _RAND_3968[31:0];
  _RAND_3969 = {1{`RANDOM}};
  reg_csr_3969 = _RAND_3969[31:0];
  _RAND_3970 = {1{`RANDOM}};
  reg_csr_3970 = _RAND_3970[31:0];
  _RAND_3971 = {1{`RANDOM}};
  reg_csr_3971 = _RAND_3971[31:0];
  _RAND_3972 = {1{`RANDOM}};
  reg_csr_3972 = _RAND_3972[31:0];
  _RAND_3973 = {1{`RANDOM}};
  reg_csr_3973 = _RAND_3973[31:0];
  _RAND_3974 = {1{`RANDOM}};
  reg_csr_3974 = _RAND_3974[31:0];
  _RAND_3975 = {1{`RANDOM}};
  reg_csr_3975 = _RAND_3975[31:0];
  _RAND_3976 = {1{`RANDOM}};
  reg_csr_3976 = _RAND_3976[31:0];
  _RAND_3977 = {1{`RANDOM}};
  reg_csr_3977 = _RAND_3977[31:0];
  _RAND_3978 = {1{`RANDOM}};
  reg_csr_3978 = _RAND_3978[31:0];
  _RAND_3979 = {1{`RANDOM}};
  reg_csr_3979 = _RAND_3979[31:0];
  _RAND_3980 = {1{`RANDOM}};
  reg_csr_3980 = _RAND_3980[31:0];
  _RAND_3981 = {1{`RANDOM}};
  reg_csr_3981 = _RAND_3981[31:0];
  _RAND_3982 = {1{`RANDOM}};
  reg_csr_3982 = _RAND_3982[31:0];
  _RAND_3983 = {1{`RANDOM}};
  reg_csr_3983 = _RAND_3983[31:0];
  _RAND_3984 = {1{`RANDOM}};
  reg_csr_3984 = _RAND_3984[31:0];
  _RAND_3985 = {1{`RANDOM}};
  reg_csr_3985 = _RAND_3985[31:0];
  _RAND_3986 = {1{`RANDOM}};
  reg_csr_3986 = _RAND_3986[31:0];
  _RAND_3987 = {1{`RANDOM}};
  reg_csr_3987 = _RAND_3987[31:0];
  _RAND_3988 = {1{`RANDOM}};
  reg_csr_3988 = _RAND_3988[31:0];
  _RAND_3989 = {1{`RANDOM}};
  reg_csr_3989 = _RAND_3989[31:0];
  _RAND_3990 = {1{`RANDOM}};
  reg_csr_3990 = _RAND_3990[31:0];
  _RAND_3991 = {1{`RANDOM}};
  reg_csr_3991 = _RAND_3991[31:0];
  _RAND_3992 = {1{`RANDOM}};
  reg_csr_3992 = _RAND_3992[31:0];
  _RAND_3993 = {1{`RANDOM}};
  reg_csr_3993 = _RAND_3993[31:0];
  _RAND_3994 = {1{`RANDOM}};
  reg_csr_3994 = _RAND_3994[31:0];
  _RAND_3995 = {1{`RANDOM}};
  reg_csr_3995 = _RAND_3995[31:0];
  _RAND_3996 = {1{`RANDOM}};
  reg_csr_3996 = _RAND_3996[31:0];
  _RAND_3997 = {1{`RANDOM}};
  reg_csr_3997 = _RAND_3997[31:0];
  _RAND_3998 = {1{`RANDOM}};
  reg_csr_3998 = _RAND_3998[31:0];
  _RAND_3999 = {1{`RANDOM}};
  reg_csr_3999 = _RAND_3999[31:0];
  _RAND_4000 = {1{`RANDOM}};
  reg_csr_4000 = _RAND_4000[31:0];
  _RAND_4001 = {1{`RANDOM}};
  reg_csr_4001 = _RAND_4001[31:0];
  _RAND_4002 = {1{`RANDOM}};
  reg_csr_4002 = _RAND_4002[31:0];
  _RAND_4003 = {1{`RANDOM}};
  reg_csr_4003 = _RAND_4003[31:0];
  _RAND_4004 = {1{`RANDOM}};
  reg_csr_4004 = _RAND_4004[31:0];
  _RAND_4005 = {1{`RANDOM}};
  reg_csr_4005 = _RAND_4005[31:0];
  _RAND_4006 = {1{`RANDOM}};
  reg_csr_4006 = _RAND_4006[31:0];
  _RAND_4007 = {1{`RANDOM}};
  reg_csr_4007 = _RAND_4007[31:0];
  _RAND_4008 = {1{`RANDOM}};
  reg_csr_4008 = _RAND_4008[31:0];
  _RAND_4009 = {1{`RANDOM}};
  reg_csr_4009 = _RAND_4009[31:0];
  _RAND_4010 = {1{`RANDOM}};
  reg_csr_4010 = _RAND_4010[31:0];
  _RAND_4011 = {1{`RANDOM}};
  reg_csr_4011 = _RAND_4011[31:0];
  _RAND_4012 = {1{`RANDOM}};
  reg_csr_4012 = _RAND_4012[31:0];
  _RAND_4013 = {1{`RANDOM}};
  reg_csr_4013 = _RAND_4013[31:0];
  _RAND_4014 = {1{`RANDOM}};
  reg_csr_4014 = _RAND_4014[31:0];
  _RAND_4015 = {1{`RANDOM}};
  reg_csr_4015 = _RAND_4015[31:0];
  _RAND_4016 = {1{`RANDOM}};
  reg_csr_4016 = _RAND_4016[31:0];
  _RAND_4017 = {1{`RANDOM}};
  reg_csr_4017 = _RAND_4017[31:0];
  _RAND_4018 = {1{`RANDOM}};
  reg_csr_4018 = _RAND_4018[31:0];
  _RAND_4019 = {1{`RANDOM}};
  reg_csr_4019 = _RAND_4019[31:0];
  _RAND_4020 = {1{`RANDOM}};
  reg_csr_4020 = _RAND_4020[31:0];
  _RAND_4021 = {1{`RANDOM}};
  reg_csr_4021 = _RAND_4021[31:0];
  _RAND_4022 = {1{`RANDOM}};
  reg_csr_4022 = _RAND_4022[31:0];
  _RAND_4023 = {1{`RANDOM}};
  reg_csr_4023 = _RAND_4023[31:0];
  _RAND_4024 = {1{`RANDOM}};
  reg_csr_4024 = _RAND_4024[31:0];
  _RAND_4025 = {1{`RANDOM}};
  reg_csr_4025 = _RAND_4025[31:0];
  _RAND_4026 = {1{`RANDOM}};
  reg_csr_4026 = _RAND_4026[31:0];
  _RAND_4027 = {1{`RANDOM}};
  reg_csr_4027 = _RAND_4027[31:0];
  _RAND_4028 = {1{`RANDOM}};
  reg_csr_4028 = _RAND_4028[31:0];
  _RAND_4029 = {1{`RANDOM}};
  reg_csr_4029 = _RAND_4029[31:0];
  _RAND_4030 = {1{`RANDOM}};
  reg_csr_4030 = _RAND_4030[31:0];
  _RAND_4031 = {1{`RANDOM}};
  reg_csr_4031 = _RAND_4031[31:0];
  _RAND_4032 = {1{`RANDOM}};
  reg_csr_4032 = _RAND_4032[31:0];
  _RAND_4033 = {1{`RANDOM}};
  reg_csr_4033 = _RAND_4033[31:0];
  _RAND_4034 = {1{`RANDOM}};
  reg_csr_4034 = _RAND_4034[31:0];
  _RAND_4035 = {1{`RANDOM}};
  reg_csr_4035 = _RAND_4035[31:0];
  _RAND_4036 = {1{`RANDOM}};
  reg_csr_4036 = _RAND_4036[31:0];
  _RAND_4037 = {1{`RANDOM}};
  reg_csr_4037 = _RAND_4037[31:0];
  _RAND_4038 = {1{`RANDOM}};
  reg_csr_4038 = _RAND_4038[31:0];
  _RAND_4039 = {1{`RANDOM}};
  reg_csr_4039 = _RAND_4039[31:0];
  _RAND_4040 = {1{`RANDOM}};
  reg_csr_4040 = _RAND_4040[31:0];
  _RAND_4041 = {1{`RANDOM}};
  reg_csr_4041 = _RAND_4041[31:0];
  _RAND_4042 = {1{`RANDOM}};
  reg_csr_4042 = _RAND_4042[31:0];
  _RAND_4043 = {1{`RANDOM}};
  reg_csr_4043 = _RAND_4043[31:0];
  _RAND_4044 = {1{`RANDOM}};
  reg_csr_4044 = _RAND_4044[31:0];
  _RAND_4045 = {1{`RANDOM}};
  reg_csr_4045 = _RAND_4045[31:0];
  _RAND_4046 = {1{`RANDOM}};
  reg_csr_4046 = _RAND_4046[31:0];
  _RAND_4047 = {1{`RANDOM}};
  reg_csr_4047 = _RAND_4047[31:0];
  _RAND_4048 = {1{`RANDOM}};
  reg_csr_4048 = _RAND_4048[31:0];
  _RAND_4049 = {1{`RANDOM}};
  reg_csr_4049 = _RAND_4049[31:0];
  _RAND_4050 = {1{`RANDOM}};
  reg_csr_4050 = _RAND_4050[31:0];
  _RAND_4051 = {1{`RANDOM}};
  reg_csr_4051 = _RAND_4051[31:0];
  _RAND_4052 = {1{`RANDOM}};
  reg_csr_4052 = _RAND_4052[31:0];
  _RAND_4053 = {1{`RANDOM}};
  reg_csr_4053 = _RAND_4053[31:0];
  _RAND_4054 = {1{`RANDOM}};
  reg_csr_4054 = _RAND_4054[31:0];
  _RAND_4055 = {1{`RANDOM}};
  reg_csr_4055 = _RAND_4055[31:0];
  _RAND_4056 = {1{`RANDOM}};
  reg_csr_4056 = _RAND_4056[31:0];
  _RAND_4057 = {1{`RANDOM}};
  reg_csr_4057 = _RAND_4057[31:0];
  _RAND_4058 = {1{`RANDOM}};
  reg_csr_4058 = _RAND_4058[31:0];
  _RAND_4059 = {1{`RANDOM}};
  reg_csr_4059 = _RAND_4059[31:0];
  _RAND_4060 = {1{`RANDOM}};
  reg_csr_4060 = _RAND_4060[31:0];
  _RAND_4061 = {1{`RANDOM}};
  reg_csr_4061 = _RAND_4061[31:0];
  _RAND_4062 = {1{`RANDOM}};
  reg_csr_4062 = _RAND_4062[31:0];
  _RAND_4063 = {1{`RANDOM}};
  reg_csr_4063 = _RAND_4063[31:0];
  _RAND_4064 = {1{`RANDOM}};
  reg_csr_4064 = _RAND_4064[31:0];
  _RAND_4065 = {1{`RANDOM}};
  reg_csr_4065 = _RAND_4065[31:0];
  _RAND_4066 = {1{`RANDOM}};
  reg_csr_4066 = _RAND_4066[31:0];
  _RAND_4067 = {1{`RANDOM}};
  reg_csr_4067 = _RAND_4067[31:0];
  _RAND_4068 = {1{`RANDOM}};
  reg_csr_4068 = _RAND_4068[31:0];
  _RAND_4069 = {1{`RANDOM}};
  reg_csr_4069 = _RAND_4069[31:0];
  _RAND_4070 = {1{`RANDOM}};
  reg_csr_4070 = _RAND_4070[31:0];
  _RAND_4071 = {1{`RANDOM}};
  reg_csr_4071 = _RAND_4071[31:0];
  _RAND_4072 = {1{`RANDOM}};
  reg_csr_4072 = _RAND_4072[31:0];
  _RAND_4073 = {1{`RANDOM}};
  reg_csr_4073 = _RAND_4073[31:0];
  _RAND_4074 = {1{`RANDOM}};
  reg_csr_4074 = _RAND_4074[31:0];
  _RAND_4075 = {1{`RANDOM}};
  reg_csr_4075 = _RAND_4075[31:0];
  _RAND_4076 = {1{`RANDOM}};
  reg_csr_4076 = _RAND_4076[31:0];
  _RAND_4077 = {1{`RANDOM}};
  reg_csr_4077 = _RAND_4077[31:0];
  _RAND_4078 = {1{`RANDOM}};
  reg_csr_4078 = _RAND_4078[31:0];
  _RAND_4079 = {1{`RANDOM}};
  reg_csr_4079 = _RAND_4079[31:0];
  _RAND_4080 = {1{`RANDOM}};
  reg_csr_4080 = _RAND_4080[31:0];
  _RAND_4081 = {1{`RANDOM}};
  reg_csr_4081 = _RAND_4081[31:0];
  _RAND_4082 = {1{`RANDOM}};
  reg_csr_4082 = _RAND_4082[31:0];
  _RAND_4083 = {1{`RANDOM}};
  reg_csr_4083 = _RAND_4083[31:0];
  _RAND_4084 = {1{`RANDOM}};
  reg_csr_4084 = _RAND_4084[31:0];
  _RAND_4085 = {1{`RANDOM}};
  reg_csr_4085 = _RAND_4085[31:0];
  _RAND_4086 = {1{`RANDOM}};
  reg_csr_4086 = _RAND_4086[31:0];
  _RAND_4087 = {1{`RANDOM}};
  reg_csr_4087 = _RAND_4087[31:0];
  _RAND_4088 = {1{`RANDOM}};
  reg_csr_4088 = _RAND_4088[31:0];
  _RAND_4089 = {1{`RANDOM}};
  reg_csr_4089 = _RAND_4089[31:0];
  _RAND_4090 = {1{`RANDOM}};
  reg_csr_4090 = _RAND_4090[31:0];
  _RAND_4091 = {1{`RANDOM}};
  reg_csr_4091 = _RAND_4091[31:0];
  _RAND_4092 = {1{`RANDOM}};
  reg_csr_4092 = _RAND_4092[31:0];
  _RAND_4093 = {1{`RANDOM}};
  reg_csr_4093 = _RAND_4093[31:0];
  _RAND_4094 = {1{`RANDOM}};
  reg_csr_4094 = _RAND_4094[31:0];
  _RAND_4095 = {1{`RANDOM}};
  reg_csr_4095 = _RAND_4095[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BR(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_io_reg_pc,
  input  [31:0] io_in_id_io_op1_data,
  input  [31:0] io_in_id_io_op2_data,
  input  [4:0]  io_in_id_io_exe_fun,
  input  [31:0] io_in_id_io_imm_b_sext,
  output        io_out_br_flag,
  output [31:0] io_out_br_target,
  output        io_out_pt_flag
);
  wire [31:0] br_target = io_in_if_io_reg_pc + io_in_id_io_imm_b_sext; // @[BR.scala 56:30]
  wire  _br_flag_T = io_in_id_io_exe_fun == 5'hb; // @[BR.scala 58:18]
  wire  _br_flag_T_1 = io_in_id_io_op1_data == io_in_id_io_op2_data; // @[BR.scala 58:45]
  wire  _br_flag_T_2 = io_in_id_io_exe_fun == 5'hc; // @[BR.scala 59:18]
  wire  _br_flag_T_4 = ~_br_flag_T_1; // @[BR.scala 59:34]
  wire  _br_flag_T_5 = io_in_id_io_exe_fun == 5'hd; // @[BR.scala 60:18]
  wire  _br_flag_T_8 = $signed(io_in_id_io_op1_data) < $signed(io_in_id_io_op2_data); // @[BR.scala 60:54]
  wire  _br_flag_T_9 = io_in_id_io_exe_fun == 5'he; // @[BR.scala 61:18]
  wire  _br_flag_T_13 = ~_br_flag_T_8; // @[BR.scala 61:34]
  wire  _br_flag_T_14 = io_in_id_io_exe_fun == 5'hf; // @[BR.scala 62:18]
  wire  _br_flag_T_15 = io_in_id_io_op1_data < io_in_id_io_op2_data; // @[BR.scala 62:45]
  wire  _br_flag_T_16 = io_in_id_io_exe_fun == 5'h10; // @[BR.scala 63:18]
  wire  _br_flag_T_18 = ~_br_flag_T_15; // @[BR.scala 63:34]
  wire  _br_flag_T_20 = _br_flag_T_14 ? _br_flag_T_15 : _br_flag_T_16 & _br_flag_T_18; // @[Mux.scala 98:16]
  wire  _br_flag_T_21 = _br_flag_T_9 ? _br_flag_T_13 : _br_flag_T_20; // @[Mux.scala 98:16]
  wire  _br_flag_T_22 = _br_flag_T_5 ? _br_flag_T_8 : _br_flag_T_21; // @[Mux.scala 98:16]
  wire  _br_flag_T_23 = _br_flag_T_2 ? _br_flag_T_4 : _br_flag_T_22; // @[Mux.scala 98:16]
  wire  br_flag = _br_flag_T ? _br_flag_T_1 : _br_flag_T_23; // @[Mux.scala 98:16]
  wire  _T_1 = ~reset; // @[BR.scala 82:11]
  assign io_out_br_flag = _br_flag_T ? _br_flag_T_1 : _br_flag_T_23; // @[Mux.scala 98:16]
  assign io_out_br_target = io_in_if_io_reg_pc + io_in_id_io_imm_b_sext; // @[BR.scala 56:30]
  assign io_out_pt_flag = _br_flag_T | (_br_flag_T_2 | (_br_flag_T_5 | (_br_flag_T_9 | (_br_flag_T_14 | _br_flag_T_16)))
    ); // @[Mux.scala 98:16]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"branch_flg: %d\n",br_flag); // @[BR.scala 82:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"branch_target: 0x%x\n",br_target); // @[BR.scala 83:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EX(
  input         clock,
  input         reset,
  input  [31:0] io_in_if_io_reg_pc,
  input  [31:0] io_in_id_io_op1_data,
  input  [31:0] io_in_id_io_op2_data,
  input  [31:0] io_in_id_io_csr_addr_default,
  input  [4:0]  io_in_id_io_exe_fun,
  input  [2:0]  io_in_id_io_rd_sel,
  input  [2:0]  io_in_id_io_csr_cmd,
  input  [31:0] io_in_id_io_imm_b_sext,
  output [31:0] io_out_alu_io_alu_out,
  output        io_out_alu_io_jump_flag,
  output [31:0] io_out_csr_io_csr_rdata,
  output [31:0] io_out_csr_io_trap_vector,
  output        io_out_br_io_br_flag,
  output [31:0] io_out_br_io_br_target,
  output        io_out_br_io_pt_flag
);
  wire  alu_clock; // @[EX.scala 46:21]
  wire  alu_reset; // @[EX.scala 46:21]
  wire [31:0] alu_io_in_id_io_op1_data; // @[EX.scala 46:21]
  wire [31:0] alu_io_in_id_io_op2_data; // @[EX.scala 46:21]
  wire [4:0] alu_io_in_id_io_exe_fun; // @[EX.scala 46:21]
  wire [2:0] alu_io_in_id_io_rd_sel; // @[EX.scala 46:21]
  wire [31:0] alu_io_out_alu_out; // @[EX.scala 46:21]
  wire  alu_io_out_jump_flag; // @[EX.scala 46:21]
  wire  csr_clock; // @[EX.scala 47:21]
  wire  csr_reset; // @[EX.scala 47:21]
  wire [31:0] csr_io_in_id_io_op1_data; // @[EX.scala 47:21]
  wire [31:0] csr_io_in_id_io_csr_addr_default; // @[EX.scala 47:21]
  wire [2:0] csr_io_in_id_io_csr_cmd; // @[EX.scala 47:21]
  wire [31:0] csr_io_out_csr_rdata; // @[EX.scala 47:21]
  wire [31:0] csr_io_out_trap_vector; // @[EX.scala 47:21]
  wire  br_clock; // @[EX.scala 48:21]
  wire  br_reset; // @[EX.scala 48:21]
  wire [31:0] br_io_in_if_io_reg_pc; // @[EX.scala 48:21]
  wire [31:0] br_io_in_id_io_op1_data; // @[EX.scala 48:21]
  wire [31:0] br_io_in_id_io_op2_data; // @[EX.scala 48:21]
  wire [4:0] br_io_in_id_io_exe_fun; // @[EX.scala 48:21]
  wire [31:0] br_io_in_id_io_imm_b_sext; // @[EX.scala 48:21]
  wire  br_io_out_br_flag; // @[EX.scala 48:21]
  wire [31:0] br_io_out_br_target; // @[EX.scala 48:21]
  wire  br_io_out_pt_flag; // @[EX.scala 48:21]
  ALU alu ( // @[EX.scala 46:21]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_id_io_op1_data(alu_io_in_id_io_op1_data),
    .io_in_id_io_op2_data(alu_io_in_id_io_op2_data),
    .io_in_id_io_exe_fun(alu_io_in_id_io_exe_fun),
    .io_in_id_io_rd_sel(alu_io_in_id_io_rd_sel),
    .io_out_alu_out(alu_io_out_alu_out),
    .io_out_jump_flag(alu_io_out_jump_flag)
  );
  CSR csr ( // @[EX.scala 47:21]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_id_io_op1_data(csr_io_in_id_io_op1_data),
    .io_in_id_io_csr_addr_default(csr_io_in_id_io_csr_addr_default),
    .io_in_id_io_csr_cmd(csr_io_in_id_io_csr_cmd),
    .io_out_csr_rdata(csr_io_out_csr_rdata),
    .io_out_trap_vector(csr_io_out_trap_vector)
  );
  BR br ( // @[EX.scala 48:21]
    .clock(br_clock),
    .reset(br_reset),
    .io_in_if_io_reg_pc(br_io_in_if_io_reg_pc),
    .io_in_id_io_op1_data(br_io_in_id_io_op1_data),
    .io_in_id_io_op2_data(br_io_in_id_io_op2_data),
    .io_in_id_io_exe_fun(br_io_in_id_io_exe_fun),
    .io_in_id_io_imm_b_sext(br_io_in_id_io_imm_b_sext),
    .io_out_br_flag(br_io_out_br_flag),
    .io_out_br_target(br_io_out_br_target),
    .io_out_pt_flag(br_io_out_pt_flag)
  );
  assign io_out_alu_io_alu_out = alu_io_out_alu_out; // @[EX.scala 59:19]
  assign io_out_alu_io_jump_flag = alu_io_out_jump_flag; // @[EX.scala 59:19]
  assign io_out_csr_io_csr_rdata = csr_io_out_csr_rdata; // @[EX.scala 60:19]
  assign io_out_csr_io_trap_vector = csr_io_out_trap_vector; // @[EX.scala 60:19]
  assign io_out_br_io_br_flag = br_io_out_br_flag; // @[EX.scala 61:19]
  assign io_out_br_io_br_target = br_io_out_br_target; // @[EX.scala 61:19]
  assign io_out_br_io_pt_flag = br_io_out_pt_flag; // @[EX.scala 61:19]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_id_io_op1_data = io_in_id_io_op1_data; // @[EX.scala 53:21]
  assign alu_io_in_id_io_op2_data = io_in_id_io_op2_data; // @[EX.scala 53:21]
  assign alu_io_in_id_io_exe_fun = io_in_id_io_exe_fun; // @[EX.scala 53:21]
  assign alu_io_in_id_io_rd_sel = io_in_id_io_rd_sel; // @[EX.scala 53:21]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_id_io_op1_data = io_in_id_io_op1_data; // @[EX.scala 54:21]
  assign csr_io_in_id_io_csr_addr_default = io_in_id_io_csr_addr_default; // @[EX.scala 54:21]
  assign csr_io_in_id_io_csr_cmd = io_in_id_io_csr_cmd; // @[EX.scala 54:21]
  assign br_clock = clock;
  assign br_reset = reset;
  assign br_io_in_if_io_reg_pc = io_in_if_io_reg_pc; // @[EX.scala 55:20]
  assign br_io_in_id_io_op1_data = io_in_id_io_op1_data; // @[EX.scala 56:20]
  assign br_io_in_id_io_op2_data = io_in_id_io_op2_data; // @[EX.scala 56:20]
  assign br_io_in_id_io_exe_fun = io_in_id_io_exe_fun; // @[EX.scala 56:20]
  assign br_io_in_id_io_imm_b_sext = io_in_id_io_imm_b_sext; // @[EX.scala 56:20]
endmodule
module MEM(
  input  [31:0] io_in_if_io_reg_pc,
  input  [4:0]  io_in_id_io_rd_addr,
  input         io_in_id_io_mem_wen,
  input         io_in_id_io_rd_wen,
  input  [2:0]  io_in_id_io_rd_sel,
  input  [31:0] io_in_id_io_rs2_data,
  input  [31:0] io_in_ex_io_alu_io_alu_out,
  input  [31:0] io_in_ex_io_csr_io_csr_rdata,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data,
  output [31:0] io_mmu_addr,
  input  [31:0] io_mmu_rdata,
  output        io_mmu_wen,
  output [31:0] io_mmu_wdata
);
  wire  _rd_data_T = io_in_id_io_rd_sel == 3'h1; // @[MEM.scala 67:17]
  wire  _rd_data_T_1 = io_in_id_io_rd_sel == 3'h2; // @[MEM.scala 68:17]
  wire [31:0] _rd_data_T_3 = io_in_if_io_reg_pc + 32'h4; // @[MEM.scala 68:40]
  wire  _rd_data_T_4 = io_in_id_io_rd_sel == 3'h3; // @[MEM.scala 69:17]
  wire [31:0] _rd_data_T_5 = _rd_data_T_4 ? io_in_ex_io_csr_io_csr_rdata : io_in_ex_io_alu_io_alu_out; // @[Mux.scala 98:16]
  wire [31:0] _rd_data_T_6 = _rd_data_T_1 ? _rd_data_T_3 : _rd_data_T_5; // @[Mux.scala 98:16]
  assign io_out_rd_wen = io_in_id_io_rd_wen; // @[MEM.scala 73:21]
  assign io_out_rd_addr = io_in_id_io_rd_addr; // @[MEM.scala 74:21]
  assign io_out_rd_data = _rd_data_T ? io_mmu_rdata : _rd_data_T_6; // @[Mux.scala 98:16]
  assign io_mmu_addr = io_in_ex_io_alu_io_alu_out; // @[MEM.scala 78:21]
  assign io_mmu_wen = io_in_id_io_mem_wen; // @[MEM.scala 77:38]
  assign io_mmu_wdata = io_in_id_io_rs2_data; // @[MEM.scala 79:21]
endmodule
module MMU(
  input  [31:0] io_mem_io_addr,
  output [31:0] io_mem_io_rdata,
  input         io_mem_io_wen,
  input  [31:0] io_mem_io_wdata,
  output [31:0] io_datamem_addr,
  input  [31:0] io_datamem_rdata,
  output        io_datamem_wen,
  output [31:0] io_datamem_wdata,
  output [31:0] io_out_apb_bus_addr,
  output        io_out_apb_bus_wen,
  output [31:0] io_out_apb_bus_wdata,
  input         io_out_apb_bus_valid,
  input  [31:0] io_out_apb_bus_rdata
);
  wire [31:0] _GEN_0 = io_out_apb_bus_valid ? io_out_apb_bus_rdata : 32'h0; // @[MMU.scala 50:25 MMU.scala 51:21 MMU.scala 53:21]
  wire  _GEN_2 = io_mem_io_addr >= 32'h10000 & io_mem_io_addr < 32'h20000 & io_mem_io_wen; // @[MMU.scala 46:84 MMU.scala 49:21 MMU.scala 58:21]
  wire [31:0] _GEN_3 = io_mem_io_addr >= 32'h10000 & io_mem_io_addr < 32'h20000 ? _GEN_0 : 32'h0; // @[MMU.scala 46:84 MMU.scala 59:21]
  assign io_mem_io_rdata = io_mem_io_addr < 32'h10000 ? io_datamem_rdata : _GEN_3; // @[MMU.scala 41:63 MMU.scala 45:21]
  assign io_datamem_addr = io_mem_io_addr - 32'h0; // @[MMU.scala 30:32]
  assign io_datamem_wen = io_mem_io_addr < 32'h10000 & io_mem_io_wen; // @[MMU.scala 41:63 MMU.scala 43:21]
  assign io_datamem_wdata = io_mem_io_wdata; // @[MMU.scala 65:25]
  assign io_out_apb_bus_addr = io_mem_io_addr - 32'h10000; // @[MMU.scala 34:25]
  assign io_out_apb_bus_wen = io_mem_io_addr < 32'h10000 ? 1'h0 : _GEN_2; // @[MMU.scala 41:63 MMU.scala 44:21]
  assign io_out_apb_bus_wdata = io_mem_io_wdata; // @[MMU.scala 69:26]
endmodule
module WB(
  input         clock,
  input         reset,
  input         io_in_mem_io_rd_wen,
  input  [4:0]  io_in_mem_io_rd_addr,
  input  [31:0] io_in_mem_io_rd_data,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data
);
  wire  _T_1 = ~reset; // @[WB.scala 60:11]
  assign io_out_rd_wen = io_in_mem_io_rd_wen; // @[WB.scala 55:21]
  assign io_out_rd_addr = io_in_mem_io_rd_addr; // @[WB.scala 56:21]
  assign io_out_rd_data = io_in_mem_io_rd_data; // @[WB.scala 57:21]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"-------------WB------------\n"); // @[WB.scala 60:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_wen: %d\n",io_in_mem_io_rd_wen); // @[WB.scala 61:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_addr: %d\n",io_in_mem_io_rd_addr); // @[WB.scala 62:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"rd_data: 0x%x\n",io_in_mem_io_rd_data); // @[WB.scala 63:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PC_BUBBLE_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_reg_pc,
  input  [31:0] io_in_inst,
  input  [31:0] io_in_ex_io_alu_io_alu_out,
  input         io_in_ex_io_alu_io_jump_flag,
  input         io_in_ex_io_br_io_br_flag,
  input  [31:0] io_in_ex_io_br_io_br_target,
  input         io_stall_io_stall_flag,
  input         io_stall_io_pred_miss_flag,
  output [31:0] io_out_reg_pc,
  output [31:0] io_out_inst,
  output [31:0] io_out_ex_io_alu_io_alu_out,
  output        io_out_ex_io_alu_io_jump_flag,
  output        io_out_ex_io_br_io_br_flag,
  output [31:0] io_out_ex_io_br_io_br_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_pc; // @[PC.scala 50:26]
  reg [31:0] inst; // @[PC.scala 51:26]
  assign io_out_reg_pc = reg_pc; // @[PC.scala 71:25]
  assign io_out_inst = inst; // @[PC.scala 72:25]
  assign io_out_ex_io_alu_io_alu_out = io_in_ex_io_alu_io_alu_out; // @[PC.scala 73:25]
  assign io_out_ex_io_alu_io_jump_flag = io_in_ex_io_alu_io_jump_flag; // @[PC.scala 73:25]
  assign io_out_ex_io_br_io_br_flag = io_in_ex_io_br_io_br_flag; // @[PC.scala 73:25]
  assign io_out_ex_io_br_io_br_target = io_in_ex_io_br_io_br_target; // @[PC.scala 73:25]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 50:26]
      reg_pc <= 32'h0; // @[PC.scala 50:26]
    end else if (!(io_stall_io_stall_flag)) begin // @[Mux.scala 98:16]
      reg_pc <= io_in_reg_pc;
    end
    if (reset) begin // @[PC.scala 51:26]
      inst <= 32'h0; // @[PC.scala 51:26]
    end else if (io_stall_io_pred_miss_flag) begin // @[Mux.scala 98:16]
      inst <= 32'h13;
    end else if (!(io_stall_io_stall_flag)) begin // @[Mux.scala 98:16]
      inst <= io_in_inst;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  inst = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PC_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_reg_pc,
  output [31:0] io_out_reg_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_io_reg_reg_pc; // @[PC.scala 30:28]
  assign io_out_reg_pc = pc_io_reg_reg_pc; // @[PC.scala 33:15]
  always @(posedge clock) begin
    if (reset) begin // @[PC.scala 30:28]
      pc_io_reg_reg_pc <= 32'h0; // @[PC.scala 30:28]
    end else begin
      pc_io_reg_reg_pc <= io_in_reg_pc; // @[PC.scala 32:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_io_reg_reg_pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ID_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_op1_data,
  input  [31:0] io_in_op2_data,
  input  [4:0]  io_in_rd_addr,
  input  [31:0] io_in_csr_addr_default,
  input  [4:0]  io_in_exe_fun,
  input         io_in_mem_wen,
  input         io_in_rd_wen,
  input  [2:0]  io_in_rd_sel,
  input  [2:0]  io_in_csr_cmd,
  input  [31:0] io_in_rs2_data,
  input  [31:0] io_in_imm_b_sext,
  output [31:0] io_out_op1_data,
  output [31:0] io_out_op2_data,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_csr_addr_default,
  output [4:0]  io_out_exe_fun,
  output        io_out_mem_wen,
  output        io_out_rd_wen,
  output [2:0]  io_out_rd_sel,
  output [2:0]  io_out_csr_cmd,
  output [31:0] io_out_rs2_data,
  output [31:0] io_out_imm_b_sext
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] id_io_reg_op1_data; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_op2_data; // @[ID.scala 53:28]
  reg [4:0] id_io_reg_rd_addr; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_csr_addr_default; // @[ID.scala 53:28]
  reg [4:0] id_io_reg_exe_fun; // @[ID.scala 53:28]
  reg  id_io_reg_mem_wen; // @[ID.scala 53:28]
  reg  id_io_reg_rd_wen; // @[ID.scala 53:28]
  reg [2:0] id_io_reg_rd_sel; // @[ID.scala 53:28]
  reg [2:0] id_io_reg_csr_cmd; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_rs2_data; // @[ID.scala 53:28]
  reg [31:0] id_io_reg_imm_b_sext; // @[ID.scala 53:28]
  assign io_out_op1_data = id_io_reg_op1_data; // @[ID.scala 56:17]
  assign io_out_op2_data = id_io_reg_op2_data; // @[ID.scala 56:17]
  assign io_out_rd_addr = id_io_reg_rd_addr; // @[ID.scala 56:17]
  assign io_out_csr_addr_default = id_io_reg_csr_addr_default; // @[ID.scala 56:17]
  assign io_out_exe_fun = id_io_reg_exe_fun; // @[ID.scala 56:17]
  assign io_out_mem_wen = id_io_reg_mem_wen; // @[ID.scala 56:17]
  assign io_out_rd_wen = id_io_reg_rd_wen; // @[ID.scala 56:17]
  assign io_out_rd_sel = id_io_reg_rd_sel; // @[ID.scala 56:17]
  assign io_out_csr_cmd = id_io_reg_csr_cmd; // @[ID.scala 56:17]
  assign io_out_rs2_data = id_io_reg_rs2_data; // @[ID.scala 56:17]
  assign io_out_imm_b_sext = id_io_reg_imm_b_sext; // @[ID.scala 56:17]
  always @(posedge clock) begin
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_op1_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_op1_data <= io_in_op1_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_op2_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_op2_data <= io_in_op2_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_addr <= 5'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_addr <= io_in_rd_addr; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_csr_addr_default <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_csr_addr_default <= io_in_csr_addr_default; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_exe_fun <= 5'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_exe_fun <= io_in_exe_fun; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_mem_wen <= 1'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_mem_wen <= io_in_mem_wen; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_wen <= 1'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_wen <= io_in_rd_wen; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rd_sel <= 3'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rd_sel <= io_in_rd_sel; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_csr_cmd <= 3'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_csr_cmd <= io_in_csr_cmd; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_rs2_data <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_rs2_data <= io_in_rs2_data; // @[ID.scala 55:17]
    end
    if (reset) begin // @[ID.scala 53:28]
      id_io_reg_imm_b_sext <= 32'h0; // @[ID.scala 53:28]
    end else begin
      id_io_reg_imm_b_sext <= io_in_imm_b_sext; // @[ID.scala 55:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  id_io_reg_op1_data = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  id_io_reg_op2_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_io_reg_rd_addr = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  id_io_reg_csr_addr_default = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  id_io_reg_exe_fun = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  id_io_reg_mem_wen = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  id_io_reg_rd_wen = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  id_io_reg_rd_sel = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  id_io_reg_csr_cmd = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  id_io_reg_rs2_data = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  id_io_reg_imm_b_sext = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EX_IO_REG(
  input         clock,
  input         reset,
  input  [31:0] io_in_alu_io_alu_out,
  input  [31:0] io_in_csr_io_csr_rdata,
  output [31:0] io_out_alu_io_alu_out,
  output [31:0] io_out_csr_io_csr_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ex_io_reg_alu_io_alu_out; // @[EX.scala 29:28]
  reg [31:0] ex_io_reg_csr_io_csr_rdata; // @[EX.scala 29:28]
  assign io_out_alu_io_alu_out = ex_io_reg_alu_io_alu_out; // @[EX.scala 32:12]
  assign io_out_csr_io_csr_rdata = ex_io_reg_csr_io_csr_rdata; // @[EX.scala 32:12]
  always @(posedge clock) begin
    if (reset) begin // @[EX.scala 29:28]
      ex_io_reg_alu_io_alu_out <= 32'h0; // @[EX.scala 29:28]
    end else begin
      ex_io_reg_alu_io_alu_out <= io_in_alu_io_alu_out; // @[EX.scala 31:15]
    end
    if (reset) begin // @[EX.scala 29:28]
      ex_io_reg_csr_io_csr_rdata <= 32'h0; // @[EX.scala 29:28]
    end else begin
      ex_io_reg_csr_io_csr_rdata <= io_in_csr_io_csr_rdata; // @[EX.scala 31:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ex_io_reg_alu_io_alu_out = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ex_io_reg_csr_io_csr_rdata = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WB_IO_REG(
  input         clock,
  input         reset,
  input         io_in_rd_wen,
  input  [4:0]  io_in_rd_addr,
  input  [31:0] io_in_rd_data,
  output        io_out_rd_wen,
  output [4:0]  io_out_rd_addr,
  output [31:0] io_out_rd_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  wb_io_reg_rd_wen; // @[WB.scala 30:28]
  reg [4:0] wb_io_reg_rd_addr; // @[WB.scala 30:28]
  reg [31:0] wb_io_reg_rd_data; // @[WB.scala 30:28]
  assign io_out_rd_wen = wb_io_reg_rd_wen; // @[WB.scala 33:17]
  assign io_out_rd_addr = wb_io_reg_rd_addr; // @[WB.scala 33:17]
  assign io_out_rd_data = wb_io_reg_rd_data; // @[WB.scala 33:17]
  always @(posedge clock) begin
    if (reset) begin // @[WB.scala 30:28]
      wb_io_reg_rd_wen <= 1'h0; // @[WB.scala 30:28]
    end else begin
      wb_io_reg_rd_wen <= io_in_rd_wen; // @[WB.scala 32:17]
    end
    if (reset) begin // @[WB.scala 30:28]
      wb_io_reg_rd_addr <= 5'h0; // @[WB.scala 30:28]
    end else begin
      wb_io_reg_rd_addr <= io_in_rd_addr; // @[WB.scala 32:17]
    end
    if (reset) begin // @[WB.scala 30:28]
      wb_io_reg_rd_data <= 32'h0; // @[WB.scala 30:28]
    end else begin
      wb_io_reg_rd_data <= io_in_rd_data; // @[WB.scala 32:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_io_reg_rd_wen = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_io_reg_rd_addr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  wb_io_reg_rd_data = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input         clock,
  input         reset,
  output [31:0] io_bus_apb_bus_addr,
  output        io_bus_apb_bus_wen,
  output [31:0] io_bus_apb_bus_wdata,
  input         io_bus_apb_bus_valid,
  input  [31:0] io_bus_apb_bus_rdata,
  output        io_exit
);
  wire  memory_clock; // @[Top.scala 17:25]
  wire [31:0] memory_io_instmem_addr; // @[Top.scala 17:25]
  wire [31:0] memory_io_instmem_inst; // @[Top.scala 17:25]
  wire [31:0] memory_io_datamem_addr; // @[Top.scala 17:25]
  wire [31:0] memory_io_datamem_rdata; // @[Top.scala 17:25]
  wire  memory_io_datamem_wen; // @[Top.scala 17:25]
  wire [31:0] memory_io_datamem_wdata; // @[Top.scala 17:25]
  wire  pc_clock; // @[Top.scala 18:25]
  wire  pc_reset; // @[Top.scala 18:25]
  wire  pc_io_in_bp_io_pred_flag; // @[Top.scala 18:25]
  wire [31:0] pc_io_in_bp_io_pred_target; // @[Top.scala 18:25]
  wire  pc_io_in_stall_io_stall_flag; // @[Top.scala 18:25]
  wire  pc_io_in_stall_io_pred_miss_flag; // @[Top.scala 18:25]
  wire [31:0] pc_io_in_ex_io_alu_io_alu_out; // @[Top.scala 18:25]
  wire  pc_io_in_ex_io_alu_io_jump_flag; // @[Top.scala 18:25]
  wire [31:0] pc_io_in_ex_io_csr_io_trap_vector; // @[Top.scala 18:25]
  wire  pc_io_in_ex_io_br_io_br_flag; // @[Top.scala 18:25]
  wire [31:0] pc_io_in_ex_io_br_io_br_target; // @[Top.scala 18:25]
  wire [31:0] pc_io_out_reg_pc; // @[Top.scala 18:25]
  wire [31:0] pc_io_out_inst; // @[Top.scala 18:25]
  wire [31:0] pc_io_out_ex_io_alu_io_alu_out; // @[Top.scala 18:25]
  wire  pc_io_out_ex_io_alu_io_jump_flag; // @[Top.scala 18:25]
  wire  pc_io_out_ex_io_br_io_br_flag; // @[Top.scala 18:25]
  wire [31:0] pc_io_out_ex_io_br_io_br_target; // @[Top.scala 18:25]
  wire [31:0] pc_io_instmem_addr; // @[Top.scala 18:25]
  wire [31:0] pc_io_instmem_inst; // @[Top.scala 18:25]
  wire  bp_clock; // @[Top.scala 19:25]
  wire  bp_reset; // @[Top.scala 19:25]
  wire [31:0] bp_io_in_pc_io_reg_pc; // @[Top.scala 19:25]
  wire [31:0] bp_io_in_pc_io_inst; // @[Top.scala 19:25]
  wire [31:0] bp_io_in_ex_pc_io_reg_pc; // @[Top.scala 19:25]
  wire [31:0] bp_io_in_ex_io_alu_io_alu_out; // @[Top.scala 19:25]
  wire  bp_io_in_ex_io_alu_io_jump_flag; // @[Top.scala 19:25]
  wire  bp_io_in_ex_io_br_io_br_flag; // @[Top.scala 19:25]
  wire [31:0] bp_io_in_ex_io_br_io_br_target; // @[Top.scala 19:25]
  wire  bp_io_in_ex_io_br_io_pt_flag; // @[Top.scala 19:25]
  wire  bp_io_out_pred_flag; // @[Top.scala 19:25]
  wire [31:0] bp_io_out_pred_target; // @[Top.scala 19:25]
  wire  id_clock; // @[Top.scala 20:25]
  wire  id_reset; // @[Top.scala 20:25]
  wire [31:0] id_io_in_if_io_reg_pc; // @[Top.scala 20:25]
  wire [31:0] id_io_in_if_io_inst; // @[Top.scala 20:25]
  wire  id_io_in_stall_io_stall_flag; // @[Top.scala 20:25]
  wire  id_io_in_stall_io_pred_miss_flag; // @[Top.scala 20:25]
  wire  id_io_in_mem_io_rd_wen; // @[Top.scala 20:25]
  wire [4:0] id_io_in_mem_io_rd_addr; // @[Top.scala 20:25]
  wire [31:0] id_io_in_mem_io_rd_data; // @[Top.scala 20:25]
  wire  id_io_in_wb_io_rd_wen; // @[Top.scala 20:25]
  wire [4:0] id_io_in_wb_io_rd_addr; // @[Top.scala 20:25]
  wire [31:0] id_io_in_wb_io_rd_data; // @[Top.scala 20:25]
  wire [31:0] id_io_out_op1_data; // @[Top.scala 20:25]
  wire [31:0] id_io_out_op2_data; // @[Top.scala 20:25]
  wire [4:0] id_io_out_rd_addr; // @[Top.scala 20:25]
  wire [31:0] id_io_out_csr_addr_default; // @[Top.scala 20:25]
  wire [4:0] id_io_out_exe_fun; // @[Top.scala 20:25]
  wire  id_io_out_mem_wen; // @[Top.scala 20:25]
  wire  id_io_out_rd_wen; // @[Top.scala 20:25]
  wire [2:0] id_io_out_rd_sel; // @[Top.scala 20:25]
  wire [2:0] id_io_out_csr_cmd; // @[Top.scala 20:25]
  wire [31:0] id_io_out_rs2_data; // @[Top.scala 20:25]
  wire [31:0] id_io_out_imm_b_sext; // @[Top.scala 20:25]
  wire [31:0] stall_io_in_if_io_reg_pc; // @[Top.scala 21:25]
  wire [31:0] stall_io_in_if_io_inst; // @[Top.scala 21:25]
  wire [31:0] stall_io_in_if_io_ex_io_alu_io_alu_out; // @[Top.scala 21:25]
  wire  stall_io_in_if_io_ex_io_alu_io_jump_flag; // @[Top.scala 21:25]
  wire  stall_io_in_if_io_ex_io_br_io_br_flag; // @[Top.scala 21:25]
  wire [31:0] stall_io_in_if_io_ex_io_br_io_br_target; // @[Top.scala 21:25]
  wire [4:0] stall_io_in_id_reg_io_rd_addr; // @[Top.scala 21:25]
  wire  stall_io_in_id_reg_io_rd_wen; // @[Top.scala 21:25]
  wire  stall_io_out_stall_flag; // @[Top.scala 21:25]
  wire  stall_io_out_pred_miss_flag; // @[Top.scala 21:25]
  wire  ex_clock; // @[Top.scala 22:25]
  wire  ex_reset; // @[Top.scala 22:25]
  wire [31:0] ex_io_in_if_io_reg_pc; // @[Top.scala 22:25]
  wire [31:0] ex_io_in_id_io_op1_data; // @[Top.scala 22:25]
  wire [31:0] ex_io_in_id_io_op2_data; // @[Top.scala 22:25]
  wire [31:0] ex_io_in_id_io_csr_addr_default; // @[Top.scala 22:25]
  wire [4:0] ex_io_in_id_io_exe_fun; // @[Top.scala 22:25]
  wire [2:0] ex_io_in_id_io_rd_sel; // @[Top.scala 22:25]
  wire [2:0] ex_io_in_id_io_csr_cmd; // @[Top.scala 22:25]
  wire [31:0] ex_io_in_id_io_imm_b_sext; // @[Top.scala 22:25]
  wire [31:0] ex_io_out_alu_io_alu_out; // @[Top.scala 22:25]
  wire  ex_io_out_alu_io_jump_flag; // @[Top.scala 22:25]
  wire [31:0] ex_io_out_csr_io_csr_rdata; // @[Top.scala 22:25]
  wire [31:0] ex_io_out_csr_io_trap_vector; // @[Top.scala 22:25]
  wire  ex_io_out_br_io_br_flag; // @[Top.scala 22:25]
  wire [31:0] ex_io_out_br_io_br_target; // @[Top.scala 22:25]
  wire  ex_io_out_br_io_pt_flag; // @[Top.scala 22:25]
  wire [31:0] mem_io_in_if_io_reg_pc; // @[Top.scala 23:25]
  wire [4:0] mem_io_in_id_io_rd_addr; // @[Top.scala 23:25]
  wire  mem_io_in_id_io_mem_wen; // @[Top.scala 23:25]
  wire  mem_io_in_id_io_rd_wen; // @[Top.scala 23:25]
  wire [2:0] mem_io_in_id_io_rd_sel; // @[Top.scala 23:25]
  wire [31:0] mem_io_in_id_io_rs2_data; // @[Top.scala 23:25]
  wire [31:0] mem_io_in_ex_io_alu_io_alu_out; // @[Top.scala 23:25]
  wire [31:0] mem_io_in_ex_io_csr_io_csr_rdata; // @[Top.scala 23:25]
  wire  mem_io_out_rd_wen; // @[Top.scala 23:25]
  wire [4:0] mem_io_out_rd_addr; // @[Top.scala 23:25]
  wire [31:0] mem_io_out_rd_data; // @[Top.scala 23:25]
  wire [31:0] mem_io_mmu_addr; // @[Top.scala 23:25]
  wire [31:0] mem_io_mmu_rdata; // @[Top.scala 23:25]
  wire  mem_io_mmu_wen; // @[Top.scala 23:25]
  wire [31:0] mem_io_mmu_wdata; // @[Top.scala 23:25]
  wire [31:0] mmu_io_mem_io_addr; // @[Top.scala 24:25]
  wire [31:0] mmu_io_mem_io_rdata; // @[Top.scala 24:25]
  wire  mmu_io_mem_io_wen; // @[Top.scala 24:25]
  wire [31:0] mmu_io_mem_io_wdata; // @[Top.scala 24:25]
  wire [31:0] mmu_io_datamem_addr; // @[Top.scala 24:25]
  wire [31:0] mmu_io_datamem_rdata; // @[Top.scala 24:25]
  wire  mmu_io_datamem_wen; // @[Top.scala 24:25]
  wire [31:0] mmu_io_datamem_wdata; // @[Top.scala 24:25]
  wire [31:0] mmu_io_out_apb_bus_addr; // @[Top.scala 24:25]
  wire  mmu_io_out_apb_bus_wen; // @[Top.scala 24:25]
  wire [31:0] mmu_io_out_apb_bus_wdata; // @[Top.scala 24:25]
  wire  mmu_io_out_apb_bus_valid; // @[Top.scala 24:25]
  wire [31:0] mmu_io_out_apb_bus_rdata; // @[Top.scala 24:25]
  wire  wb_clock; // @[Top.scala 25:25]
  wire  wb_reset; // @[Top.scala 25:25]
  wire  wb_io_in_mem_io_rd_wen; // @[Top.scala 25:25]
  wire [4:0] wb_io_in_mem_io_rd_addr; // @[Top.scala 25:25]
  wire [31:0] wb_io_in_mem_io_rd_data; // @[Top.scala 25:25]
  wire  wb_io_out_rd_wen; // @[Top.scala 25:25]
  wire [4:0] wb_io_out_rd_addr; // @[Top.scala 25:25]
  wire [31:0] wb_io_out_rd_data; // @[Top.scala 25:25]
  wire  if_io_reg_clock; // @[Top.scala 28:33]
  wire  if_io_reg_reset; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_in_reg_pc; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_in_inst; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_in_ex_io_alu_io_alu_out; // @[Top.scala 28:33]
  wire  if_io_reg_io_in_ex_io_alu_io_jump_flag; // @[Top.scala 28:33]
  wire  if_io_reg_io_in_ex_io_br_io_br_flag; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_in_ex_io_br_io_br_target; // @[Top.scala 28:33]
  wire  if_io_reg_io_stall_io_stall_flag; // @[Top.scala 28:33]
  wire  if_io_reg_io_stall_io_pred_miss_flag; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_out_reg_pc; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_out_inst; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_out_ex_io_alu_io_alu_out; // @[Top.scala 28:33]
  wire  if_io_reg_io_out_ex_io_alu_io_jump_flag; // @[Top.scala 28:33]
  wire  if_io_reg_io_out_ex_io_br_io_br_flag; // @[Top.scala 28:33]
  wire [31:0] if_io_reg_io_out_ex_io_br_io_br_target; // @[Top.scala 28:33]
  wire  if_io_reg_n_clock; // @[Top.scala 29:33]
  wire  if_io_reg_n_reset; // @[Top.scala 29:33]
  wire [31:0] if_io_reg_n_io_in_reg_pc; // @[Top.scala 29:33]
  wire [31:0] if_io_reg_n_io_out_reg_pc; // @[Top.scala 29:33]
  wire  if_io_reg_nn_clock; // @[Top.scala 30:33]
  wire  if_io_reg_nn_reset; // @[Top.scala 30:33]
  wire [31:0] if_io_reg_nn_io_in_reg_pc; // @[Top.scala 30:33]
  wire [31:0] if_io_reg_nn_io_out_reg_pc; // @[Top.scala 30:33]
  wire  id_io_reg_clock; // @[Top.scala 31:33]
  wire  id_io_reg_reset; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_in_op1_data; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_in_op2_data; // @[Top.scala 31:33]
  wire [4:0] id_io_reg_io_in_rd_addr; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_in_csr_addr_default; // @[Top.scala 31:33]
  wire [4:0] id_io_reg_io_in_exe_fun; // @[Top.scala 31:33]
  wire  id_io_reg_io_in_mem_wen; // @[Top.scala 31:33]
  wire  id_io_reg_io_in_rd_wen; // @[Top.scala 31:33]
  wire [2:0] id_io_reg_io_in_rd_sel; // @[Top.scala 31:33]
  wire [2:0] id_io_reg_io_in_csr_cmd; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_in_rs2_data; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_in_imm_b_sext; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_out_op1_data; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_out_op2_data; // @[Top.scala 31:33]
  wire [4:0] id_io_reg_io_out_rd_addr; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_out_csr_addr_default; // @[Top.scala 31:33]
  wire [4:0] id_io_reg_io_out_exe_fun; // @[Top.scala 31:33]
  wire  id_io_reg_io_out_mem_wen; // @[Top.scala 31:33]
  wire  id_io_reg_io_out_rd_wen; // @[Top.scala 31:33]
  wire [2:0] id_io_reg_io_out_rd_sel; // @[Top.scala 31:33]
  wire [2:0] id_io_reg_io_out_csr_cmd; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_out_rs2_data; // @[Top.scala 31:33]
  wire [31:0] id_io_reg_io_out_imm_b_sext; // @[Top.scala 31:33]
  wire  id_io_reg_n_clock; // @[Top.scala 32:33]
  wire  id_io_reg_n_reset; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_in_op1_data; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_in_op2_data; // @[Top.scala 32:33]
  wire [4:0] id_io_reg_n_io_in_rd_addr; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_in_csr_addr_default; // @[Top.scala 32:33]
  wire [4:0] id_io_reg_n_io_in_exe_fun; // @[Top.scala 32:33]
  wire  id_io_reg_n_io_in_mem_wen; // @[Top.scala 32:33]
  wire  id_io_reg_n_io_in_rd_wen; // @[Top.scala 32:33]
  wire [2:0] id_io_reg_n_io_in_rd_sel; // @[Top.scala 32:33]
  wire [2:0] id_io_reg_n_io_in_csr_cmd; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_in_rs2_data; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_in_imm_b_sext; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_out_op1_data; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_out_op2_data; // @[Top.scala 32:33]
  wire [4:0] id_io_reg_n_io_out_rd_addr; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_out_csr_addr_default; // @[Top.scala 32:33]
  wire [4:0] id_io_reg_n_io_out_exe_fun; // @[Top.scala 32:33]
  wire  id_io_reg_n_io_out_mem_wen; // @[Top.scala 32:33]
  wire  id_io_reg_n_io_out_rd_wen; // @[Top.scala 32:33]
  wire [2:0] id_io_reg_n_io_out_rd_sel; // @[Top.scala 32:33]
  wire [2:0] id_io_reg_n_io_out_csr_cmd; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_out_rs2_data; // @[Top.scala 32:33]
  wire [31:0] id_io_reg_n_io_out_imm_b_sext; // @[Top.scala 32:33]
  wire  ex_io_reg_clock; // @[Top.scala 33:33]
  wire  ex_io_reg_reset; // @[Top.scala 33:33]
  wire [31:0] ex_io_reg_io_in_alu_io_alu_out; // @[Top.scala 33:33]
  wire [31:0] ex_io_reg_io_in_csr_io_csr_rdata; // @[Top.scala 33:33]
  wire [31:0] ex_io_reg_io_out_alu_io_alu_out; // @[Top.scala 33:33]
  wire [31:0] ex_io_reg_io_out_csr_io_csr_rdata; // @[Top.scala 33:33]
  wire  mem_io_reg_clock; // @[Top.scala 34:33]
  wire  mem_io_reg_reset; // @[Top.scala 34:33]
  wire  mem_io_reg_io_in_rd_wen; // @[Top.scala 34:33]
  wire [4:0] mem_io_reg_io_in_rd_addr; // @[Top.scala 34:33]
  wire [31:0] mem_io_reg_io_in_rd_data; // @[Top.scala 34:33]
  wire  mem_io_reg_io_out_rd_wen; // @[Top.scala 34:33]
  wire [4:0] mem_io_reg_io_out_rd_addr; // @[Top.scala 34:33]
  wire [31:0] mem_io_reg_io_out_rd_data; // @[Top.scala 34:33]
  wire [31:0] _io_exit_T = pc_io_out_inst; // @[Top.scala 82:17]
  wire  _io_exit_T_1 = 32'hc0001073 == _io_exit_T; // @[Top.scala 82:17]
  wire  _io_exit_T_2 = pc_io_out_inst == 32'h0; // @[Top.scala 83:17]
  wire  _io_exit_T_3 = pc_io_out_reg_pc == 32'h44; // @[Top.scala 84:17]
  Memory memory ( // @[Top.scala 17:25]
    .clock(memory_clock),
    .io_instmem_addr(memory_io_instmem_addr),
    .io_instmem_inst(memory_io_instmem_inst),
    .io_datamem_addr(memory_io_datamem_addr),
    .io_datamem_rdata(memory_io_datamem_rdata),
    .io_datamem_wen(memory_io_datamem_wen),
    .io_datamem_wdata(memory_io_datamem_wdata)
  );
  PC pc ( // @[Top.scala 18:25]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_in_bp_io_pred_flag(pc_io_in_bp_io_pred_flag),
    .io_in_bp_io_pred_target(pc_io_in_bp_io_pred_target),
    .io_in_stall_io_stall_flag(pc_io_in_stall_io_stall_flag),
    .io_in_stall_io_pred_miss_flag(pc_io_in_stall_io_pred_miss_flag),
    .io_in_ex_io_alu_io_alu_out(pc_io_in_ex_io_alu_io_alu_out),
    .io_in_ex_io_alu_io_jump_flag(pc_io_in_ex_io_alu_io_jump_flag),
    .io_in_ex_io_csr_io_trap_vector(pc_io_in_ex_io_csr_io_trap_vector),
    .io_in_ex_io_br_io_br_flag(pc_io_in_ex_io_br_io_br_flag),
    .io_in_ex_io_br_io_br_target(pc_io_in_ex_io_br_io_br_target),
    .io_out_reg_pc(pc_io_out_reg_pc),
    .io_out_inst(pc_io_out_inst),
    .io_out_ex_io_alu_io_alu_out(pc_io_out_ex_io_alu_io_alu_out),
    .io_out_ex_io_alu_io_jump_flag(pc_io_out_ex_io_alu_io_jump_flag),
    .io_out_ex_io_br_io_br_flag(pc_io_out_ex_io_br_io_br_flag),
    .io_out_ex_io_br_io_br_target(pc_io_out_ex_io_br_io_br_target),
    .io_instmem_addr(pc_io_instmem_addr),
    .io_instmem_inst(pc_io_instmem_inst)
  );
  BP bp ( // @[Top.scala 19:25]
    .clock(bp_clock),
    .reset(bp_reset),
    .io_in_pc_io_reg_pc(bp_io_in_pc_io_reg_pc),
    .io_in_pc_io_inst(bp_io_in_pc_io_inst),
    .io_in_ex_pc_io_reg_pc(bp_io_in_ex_pc_io_reg_pc),
    .io_in_ex_io_alu_io_alu_out(bp_io_in_ex_io_alu_io_alu_out),
    .io_in_ex_io_alu_io_jump_flag(bp_io_in_ex_io_alu_io_jump_flag),
    .io_in_ex_io_br_io_br_flag(bp_io_in_ex_io_br_io_br_flag),
    .io_in_ex_io_br_io_br_target(bp_io_in_ex_io_br_io_br_target),
    .io_in_ex_io_br_io_pt_flag(bp_io_in_ex_io_br_io_pt_flag),
    .io_out_pred_flag(bp_io_out_pred_flag),
    .io_out_pred_target(bp_io_out_pred_target)
  );
  ID id ( // @[Top.scala 20:25]
    .clock(id_clock),
    .reset(id_reset),
    .io_in_if_io_reg_pc(id_io_in_if_io_reg_pc),
    .io_in_if_io_inst(id_io_in_if_io_inst),
    .io_in_stall_io_stall_flag(id_io_in_stall_io_stall_flag),
    .io_in_stall_io_pred_miss_flag(id_io_in_stall_io_pred_miss_flag),
    .io_in_mem_io_rd_wen(id_io_in_mem_io_rd_wen),
    .io_in_mem_io_rd_addr(id_io_in_mem_io_rd_addr),
    .io_in_mem_io_rd_data(id_io_in_mem_io_rd_data),
    .io_in_wb_io_rd_wen(id_io_in_wb_io_rd_wen),
    .io_in_wb_io_rd_addr(id_io_in_wb_io_rd_addr),
    .io_in_wb_io_rd_data(id_io_in_wb_io_rd_data),
    .io_out_op1_data(id_io_out_op1_data),
    .io_out_op2_data(id_io_out_op2_data),
    .io_out_rd_addr(id_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_out_exe_fun),
    .io_out_mem_wen(id_io_out_mem_wen),
    .io_out_rd_wen(id_io_out_rd_wen),
    .io_out_rd_sel(id_io_out_rd_sel),
    .io_out_csr_cmd(id_io_out_csr_cmd),
    .io_out_rs2_data(id_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_out_imm_b_sext)
  );
  Stall stall ( // @[Top.scala 21:25]
    .io_in_if_io_reg_pc(stall_io_in_if_io_reg_pc),
    .io_in_if_io_inst(stall_io_in_if_io_inst),
    .io_in_if_io_ex_io_alu_io_alu_out(stall_io_in_if_io_ex_io_alu_io_alu_out),
    .io_in_if_io_ex_io_alu_io_jump_flag(stall_io_in_if_io_ex_io_alu_io_jump_flag),
    .io_in_if_io_ex_io_br_io_br_flag(stall_io_in_if_io_ex_io_br_io_br_flag),
    .io_in_if_io_ex_io_br_io_br_target(stall_io_in_if_io_ex_io_br_io_br_target),
    .io_in_id_reg_io_rd_addr(stall_io_in_id_reg_io_rd_addr),
    .io_in_id_reg_io_rd_wen(stall_io_in_id_reg_io_rd_wen),
    .io_out_stall_flag(stall_io_out_stall_flag),
    .io_out_pred_miss_flag(stall_io_out_pred_miss_flag)
  );
  EX ex ( // @[Top.scala 22:25]
    .clock(ex_clock),
    .reset(ex_reset),
    .io_in_if_io_reg_pc(ex_io_in_if_io_reg_pc),
    .io_in_id_io_op1_data(ex_io_in_id_io_op1_data),
    .io_in_id_io_op2_data(ex_io_in_id_io_op2_data),
    .io_in_id_io_csr_addr_default(ex_io_in_id_io_csr_addr_default),
    .io_in_id_io_exe_fun(ex_io_in_id_io_exe_fun),
    .io_in_id_io_rd_sel(ex_io_in_id_io_rd_sel),
    .io_in_id_io_csr_cmd(ex_io_in_id_io_csr_cmd),
    .io_in_id_io_imm_b_sext(ex_io_in_id_io_imm_b_sext),
    .io_out_alu_io_alu_out(ex_io_out_alu_io_alu_out),
    .io_out_alu_io_jump_flag(ex_io_out_alu_io_jump_flag),
    .io_out_csr_io_csr_rdata(ex_io_out_csr_io_csr_rdata),
    .io_out_csr_io_trap_vector(ex_io_out_csr_io_trap_vector),
    .io_out_br_io_br_flag(ex_io_out_br_io_br_flag),
    .io_out_br_io_br_target(ex_io_out_br_io_br_target),
    .io_out_br_io_pt_flag(ex_io_out_br_io_pt_flag)
  );
  MEM mem ( // @[Top.scala 23:25]
    .io_in_if_io_reg_pc(mem_io_in_if_io_reg_pc),
    .io_in_id_io_rd_addr(mem_io_in_id_io_rd_addr),
    .io_in_id_io_mem_wen(mem_io_in_id_io_mem_wen),
    .io_in_id_io_rd_wen(mem_io_in_id_io_rd_wen),
    .io_in_id_io_rd_sel(mem_io_in_id_io_rd_sel),
    .io_in_id_io_rs2_data(mem_io_in_id_io_rs2_data),
    .io_in_ex_io_alu_io_alu_out(mem_io_in_ex_io_alu_io_alu_out),
    .io_in_ex_io_csr_io_csr_rdata(mem_io_in_ex_io_csr_io_csr_rdata),
    .io_out_rd_wen(mem_io_out_rd_wen),
    .io_out_rd_addr(mem_io_out_rd_addr),
    .io_out_rd_data(mem_io_out_rd_data),
    .io_mmu_addr(mem_io_mmu_addr),
    .io_mmu_rdata(mem_io_mmu_rdata),
    .io_mmu_wen(mem_io_mmu_wen),
    .io_mmu_wdata(mem_io_mmu_wdata)
  );
  MMU mmu ( // @[Top.scala 24:25]
    .io_mem_io_addr(mmu_io_mem_io_addr),
    .io_mem_io_rdata(mmu_io_mem_io_rdata),
    .io_mem_io_wen(mmu_io_mem_io_wen),
    .io_mem_io_wdata(mmu_io_mem_io_wdata),
    .io_datamem_addr(mmu_io_datamem_addr),
    .io_datamem_rdata(mmu_io_datamem_rdata),
    .io_datamem_wen(mmu_io_datamem_wen),
    .io_datamem_wdata(mmu_io_datamem_wdata),
    .io_out_apb_bus_addr(mmu_io_out_apb_bus_addr),
    .io_out_apb_bus_wen(mmu_io_out_apb_bus_wen),
    .io_out_apb_bus_wdata(mmu_io_out_apb_bus_wdata),
    .io_out_apb_bus_valid(mmu_io_out_apb_bus_valid),
    .io_out_apb_bus_rdata(mmu_io_out_apb_bus_rdata)
  );
  WB wb ( // @[Top.scala 25:25]
    .clock(wb_clock),
    .reset(wb_reset),
    .io_in_mem_io_rd_wen(wb_io_in_mem_io_rd_wen),
    .io_in_mem_io_rd_addr(wb_io_in_mem_io_rd_addr),
    .io_in_mem_io_rd_data(wb_io_in_mem_io_rd_data),
    .io_out_rd_wen(wb_io_out_rd_wen),
    .io_out_rd_addr(wb_io_out_rd_addr),
    .io_out_rd_data(wb_io_out_rd_data)
  );
  PC_BUBBLE_REG if_io_reg ( // @[Top.scala 28:33]
    .clock(if_io_reg_clock),
    .reset(if_io_reg_reset),
    .io_in_reg_pc(if_io_reg_io_in_reg_pc),
    .io_in_inst(if_io_reg_io_in_inst),
    .io_in_ex_io_alu_io_alu_out(if_io_reg_io_in_ex_io_alu_io_alu_out),
    .io_in_ex_io_alu_io_jump_flag(if_io_reg_io_in_ex_io_alu_io_jump_flag),
    .io_in_ex_io_br_io_br_flag(if_io_reg_io_in_ex_io_br_io_br_flag),
    .io_in_ex_io_br_io_br_target(if_io_reg_io_in_ex_io_br_io_br_target),
    .io_stall_io_stall_flag(if_io_reg_io_stall_io_stall_flag),
    .io_stall_io_pred_miss_flag(if_io_reg_io_stall_io_pred_miss_flag),
    .io_out_reg_pc(if_io_reg_io_out_reg_pc),
    .io_out_inst(if_io_reg_io_out_inst),
    .io_out_ex_io_alu_io_alu_out(if_io_reg_io_out_ex_io_alu_io_alu_out),
    .io_out_ex_io_alu_io_jump_flag(if_io_reg_io_out_ex_io_alu_io_jump_flag),
    .io_out_ex_io_br_io_br_flag(if_io_reg_io_out_ex_io_br_io_br_flag),
    .io_out_ex_io_br_io_br_target(if_io_reg_io_out_ex_io_br_io_br_target)
  );
  PC_IO_REG if_io_reg_n ( // @[Top.scala 29:33]
    .clock(if_io_reg_n_clock),
    .reset(if_io_reg_n_reset),
    .io_in_reg_pc(if_io_reg_n_io_in_reg_pc),
    .io_out_reg_pc(if_io_reg_n_io_out_reg_pc)
  );
  PC_IO_REG if_io_reg_nn ( // @[Top.scala 30:33]
    .clock(if_io_reg_nn_clock),
    .reset(if_io_reg_nn_reset),
    .io_in_reg_pc(if_io_reg_nn_io_in_reg_pc),
    .io_out_reg_pc(if_io_reg_nn_io_out_reg_pc)
  );
  ID_IO_REG id_io_reg ( // @[Top.scala 31:33]
    .clock(id_io_reg_clock),
    .reset(id_io_reg_reset),
    .io_in_op1_data(id_io_reg_io_in_op1_data),
    .io_in_op2_data(id_io_reg_io_in_op2_data),
    .io_in_rd_addr(id_io_reg_io_in_rd_addr),
    .io_in_csr_addr_default(id_io_reg_io_in_csr_addr_default),
    .io_in_exe_fun(id_io_reg_io_in_exe_fun),
    .io_in_mem_wen(id_io_reg_io_in_mem_wen),
    .io_in_rd_wen(id_io_reg_io_in_rd_wen),
    .io_in_rd_sel(id_io_reg_io_in_rd_sel),
    .io_in_csr_cmd(id_io_reg_io_in_csr_cmd),
    .io_in_rs2_data(id_io_reg_io_in_rs2_data),
    .io_in_imm_b_sext(id_io_reg_io_in_imm_b_sext),
    .io_out_op1_data(id_io_reg_io_out_op1_data),
    .io_out_op2_data(id_io_reg_io_out_op2_data),
    .io_out_rd_addr(id_io_reg_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_reg_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_reg_io_out_exe_fun),
    .io_out_mem_wen(id_io_reg_io_out_mem_wen),
    .io_out_rd_wen(id_io_reg_io_out_rd_wen),
    .io_out_rd_sel(id_io_reg_io_out_rd_sel),
    .io_out_csr_cmd(id_io_reg_io_out_csr_cmd),
    .io_out_rs2_data(id_io_reg_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_reg_io_out_imm_b_sext)
  );
  ID_IO_REG id_io_reg_n ( // @[Top.scala 32:33]
    .clock(id_io_reg_n_clock),
    .reset(id_io_reg_n_reset),
    .io_in_op1_data(id_io_reg_n_io_in_op1_data),
    .io_in_op2_data(id_io_reg_n_io_in_op2_data),
    .io_in_rd_addr(id_io_reg_n_io_in_rd_addr),
    .io_in_csr_addr_default(id_io_reg_n_io_in_csr_addr_default),
    .io_in_exe_fun(id_io_reg_n_io_in_exe_fun),
    .io_in_mem_wen(id_io_reg_n_io_in_mem_wen),
    .io_in_rd_wen(id_io_reg_n_io_in_rd_wen),
    .io_in_rd_sel(id_io_reg_n_io_in_rd_sel),
    .io_in_csr_cmd(id_io_reg_n_io_in_csr_cmd),
    .io_in_rs2_data(id_io_reg_n_io_in_rs2_data),
    .io_in_imm_b_sext(id_io_reg_n_io_in_imm_b_sext),
    .io_out_op1_data(id_io_reg_n_io_out_op1_data),
    .io_out_op2_data(id_io_reg_n_io_out_op2_data),
    .io_out_rd_addr(id_io_reg_n_io_out_rd_addr),
    .io_out_csr_addr_default(id_io_reg_n_io_out_csr_addr_default),
    .io_out_exe_fun(id_io_reg_n_io_out_exe_fun),
    .io_out_mem_wen(id_io_reg_n_io_out_mem_wen),
    .io_out_rd_wen(id_io_reg_n_io_out_rd_wen),
    .io_out_rd_sel(id_io_reg_n_io_out_rd_sel),
    .io_out_csr_cmd(id_io_reg_n_io_out_csr_cmd),
    .io_out_rs2_data(id_io_reg_n_io_out_rs2_data),
    .io_out_imm_b_sext(id_io_reg_n_io_out_imm_b_sext)
  );
  EX_IO_REG ex_io_reg ( // @[Top.scala 33:33]
    .clock(ex_io_reg_clock),
    .reset(ex_io_reg_reset),
    .io_in_alu_io_alu_out(ex_io_reg_io_in_alu_io_alu_out),
    .io_in_csr_io_csr_rdata(ex_io_reg_io_in_csr_io_csr_rdata),
    .io_out_alu_io_alu_out(ex_io_reg_io_out_alu_io_alu_out),
    .io_out_csr_io_csr_rdata(ex_io_reg_io_out_csr_io_csr_rdata)
  );
  WB_IO_REG mem_io_reg ( // @[Top.scala 34:33]
    .clock(mem_io_reg_clock),
    .reset(mem_io_reg_reset),
    .io_in_rd_wen(mem_io_reg_io_in_rd_wen),
    .io_in_rd_addr(mem_io_reg_io_in_rd_addr),
    .io_in_rd_data(mem_io_reg_io_in_rd_data),
    .io_out_rd_wen(mem_io_reg_io_out_rd_wen),
    .io_out_rd_addr(mem_io_reg_io_out_rd_addr),
    .io_out_rd_data(mem_io_reg_io_out_rd_data)
  );
  assign io_bus_apb_bus_addr = mmu_io_out_apb_bus_addr; // @[Top.scala 86:12]
  assign io_bus_apb_bus_wen = mmu_io_out_apb_bus_wen; // @[Top.scala 86:12]
  assign io_bus_apb_bus_wdata = mmu_io_out_apb_bus_wdata; // @[Top.scala 86:12]
  assign io_exit = _io_exit_T_1 | (_io_exit_T_2 | _io_exit_T_3); // @[Mux.scala 98:16]
  assign memory_clock = clock;
  assign memory_io_instmem_addr = pc_io_instmem_addr; // @[Top.scala 40:25]
  assign memory_io_datamem_addr = mmu_io_datamem_addr; // @[Top.scala 74:25]
  assign memory_io_datamem_wen = mmu_io_datamem_wen; // @[Top.scala 74:25]
  assign memory_io_datamem_wdata = mmu_io_datamem_wdata; // @[Top.scala 74:25]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_in_bp_io_pred_flag = bp_io_out_pred_flag; // @[Top.scala 41:25]
  assign pc_io_in_bp_io_pred_target = bp_io_out_pred_target; // @[Top.scala 41:25]
  assign pc_io_in_stall_io_stall_flag = stall_io_out_stall_flag; // @[Top.scala 38:25]
  assign pc_io_in_stall_io_pred_miss_flag = stall_io_out_pred_miss_flag; // @[Top.scala 38:25]
  assign pc_io_in_ex_io_alu_io_alu_out = ex_io_out_alu_io_alu_out; // @[Top.scala 39:25]
  assign pc_io_in_ex_io_alu_io_jump_flag = ex_io_out_alu_io_jump_flag; // @[Top.scala 39:25]
  assign pc_io_in_ex_io_csr_io_trap_vector = ex_io_out_csr_io_trap_vector; // @[Top.scala 39:25]
  assign pc_io_in_ex_io_br_io_br_flag = ex_io_out_br_io_br_flag; // @[Top.scala 39:25]
  assign pc_io_in_ex_io_br_io_br_target = ex_io_out_br_io_br_target; // @[Top.scala 39:25]
  assign pc_io_instmem_inst = memory_io_instmem_inst; // @[Top.scala 40:25]
  assign bp_clock = clock;
  assign bp_reset = reset;
  assign bp_io_in_pc_io_reg_pc = pc_io_out_reg_pc; // @[Top.scala 43:25]
  assign bp_io_in_pc_io_inst = pc_io_out_inst; // @[Top.scala 43:25]
  assign bp_io_in_ex_pc_io_reg_pc = if_io_reg_n_io_out_reg_pc; // @[Top.scala 44:25]
  assign bp_io_in_ex_io_alu_io_alu_out = ex_io_out_alu_io_alu_out; // @[Top.scala 46:25]
  assign bp_io_in_ex_io_alu_io_jump_flag = ex_io_out_alu_io_jump_flag; // @[Top.scala 46:25]
  assign bp_io_in_ex_io_br_io_br_flag = ex_io_out_br_io_br_flag; // @[Top.scala 46:25]
  assign bp_io_in_ex_io_br_io_br_target = ex_io_out_br_io_br_target; // @[Top.scala 46:25]
  assign bp_io_in_ex_io_br_io_pt_flag = ex_io_out_br_io_pt_flag; // @[Top.scala 46:25]
  assign id_clock = clock;
  assign id_reset = reset;
  assign id_io_in_if_io_reg_pc = if_io_reg_io_out_reg_pc; // @[Top.scala 56:25]
  assign id_io_in_if_io_inst = if_io_reg_io_out_inst; // @[Top.scala 56:25]
  assign id_io_in_stall_io_stall_flag = stall_io_out_stall_flag; // @[Top.scala 58:25]
  assign id_io_in_stall_io_pred_miss_flag = stall_io_out_pred_miss_flag; // @[Top.scala 58:25]
  assign id_io_in_mem_io_rd_wen = mem_io_out_rd_wen; // @[Top.scala 60:25]
  assign id_io_in_mem_io_rd_addr = mem_io_out_rd_addr; // @[Top.scala 60:25]
  assign id_io_in_mem_io_rd_data = mem_io_out_rd_data; // @[Top.scala 60:25]
  assign id_io_in_wb_io_rd_wen = wb_io_out_rd_wen; // @[Top.scala 59:25]
  assign id_io_in_wb_io_rd_addr = wb_io_out_rd_addr; // @[Top.scala 59:25]
  assign id_io_in_wb_io_rd_data = wb_io_out_rd_data; // @[Top.scala 59:25]
  assign stall_io_in_if_io_reg_pc = if_io_reg_io_out_reg_pc; // @[Top.scala 49:25]
  assign stall_io_in_if_io_inst = if_io_reg_io_out_inst; // @[Top.scala 49:25]
  assign stall_io_in_if_io_ex_io_alu_io_alu_out = if_io_reg_io_out_ex_io_alu_io_alu_out; // @[Top.scala 49:25]
  assign stall_io_in_if_io_ex_io_alu_io_jump_flag = if_io_reg_io_out_ex_io_alu_io_jump_flag; // @[Top.scala 49:25]
  assign stall_io_in_if_io_ex_io_br_io_br_flag = if_io_reg_io_out_ex_io_br_io_br_flag; // @[Top.scala 49:25]
  assign stall_io_in_if_io_ex_io_br_io_br_target = if_io_reg_io_out_ex_io_br_io_br_target; // @[Top.scala 49:25]
  assign stall_io_in_id_reg_io_rd_addr = id_io_reg_io_out_rd_addr; // @[Top.scala 51:29]
  assign stall_io_in_id_reg_io_rd_wen = id_io_reg_io_out_rd_wen; // @[Top.scala 51:29]
  assign ex_clock = clock;
  assign ex_reset = reset;
  assign ex_io_in_if_io_reg_pc = if_io_reg_n_io_out_reg_pc; // @[Top.scala 64:25]
  assign ex_io_in_id_io_op1_data = id_io_reg_io_out_op1_data; // @[Top.scala 62:25]
  assign ex_io_in_id_io_op2_data = id_io_reg_io_out_op2_data; // @[Top.scala 62:25]
  assign ex_io_in_id_io_csr_addr_default = id_io_reg_io_out_csr_addr_default; // @[Top.scala 62:25]
  assign ex_io_in_id_io_exe_fun = id_io_reg_io_out_exe_fun; // @[Top.scala 62:25]
  assign ex_io_in_id_io_rd_sel = id_io_reg_io_out_rd_sel; // @[Top.scala 62:25]
  assign ex_io_in_id_io_csr_cmd = id_io_reg_io_out_csr_cmd; // @[Top.scala 62:25]
  assign ex_io_in_id_io_imm_b_sext = id_io_reg_io_out_imm_b_sext; // @[Top.scala 62:25]
  assign mem_io_in_if_io_reg_pc = if_io_reg_nn_io_out_reg_pc; // @[Top.scala 66:25]
  assign mem_io_in_id_io_rd_addr = id_io_reg_n_io_out_rd_addr; // @[Top.scala 68:25]
  assign mem_io_in_id_io_mem_wen = id_io_reg_n_io_out_mem_wen; // @[Top.scala 68:25]
  assign mem_io_in_id_io_rd_wen = id_io_reg_n_io_out_rd_wen; // @[Top.scala 68:25]
  assign mem_io_in_id_io_rd_sel = id_io_reg_n_io_out_rd_sel; // @[Top.scala 68:25]
  assign mem_io_in_id_io_rs2_data = id_io_reg_n_io_out_rs2_data; // @[Top.scala 68:25]
  assign mem_io_in_ex_io_alu_io_alu_out = ex_io_reg_io_out_alu_io_alu_out; // @[Top.scala 70:25]
  assign mem_io_in_ex_io_csr_io_csr_rdata = ex_io_reg_io_out_csr_io_csr_rdata; // @[Top.scala 70:25]
  assign mem_io_mmu_rdata = mmu_io_mem_io_rdata; // @[Top.scala 73:25]
  assign mmu_io_mem_io_addr = mem_io_mmu_addr; // @[Top.scala 73:25]
  assign mmu_io_mem_io_wen = mem_io_mmu_wen; // @[Top.scala 73:25]
  assign mmu_io_mem_io_wdata = mem_io_mmu_wdata; // @[Top.scala 73:25]
  assign mmu_io_datamem_rdata = memory_io_datamem_rdata; // @[Top.scala 74:25]
  assign mmu_io_out_apb_bus_valid = io_bus_apb_bus_valid; // @[Top.scala 86:12]
  assign mmu_io_out_apb_bus_rdata = io_bus_apb_bus_rdata; // @[Top.scala 86:12]
  assign wb_clock = clock;
  assign wb_reset = reset;
  assign wb_io_in_mem_io_rd_wen = mem_io_reg_io_out_rd_wen; // @[Top.scala 76:25]
  assign wb_io_in_mem_io_rd_addr = mem_io_reg_io_out_rd_addr; // @[Top.scala 76:25]
  assign wb_io_in_mem_io_rd_data = mem_io_reg_io_out_rd_data; // @[Top.scala 76:25]
  assign if_io_reg_clock = clock;
  assign if_io_reg_reset = reset;
  assign if_io_reg_io_in_reg_pc = pc_io_out_reg_pc; // @[Top.scala 57:29]
  assign if_io_reg_io_in_inst = pc_io_out_inst; // @[Top.scala 57:29]
  assign if_io_reg_io_in_ex_io_alu_io_alu_out = pc_io_out_ex_io_alu_io_alu_out; // @[Top.scala 57:29]
  assign if_io_reg_io_in_ex_io_alu_io_jump_flag = pc_io_out_ex_io_alu_io_jump_flag; // @[Top.scala 57:29]
  assign if_io_reg_io_in_ex_io_br_io_br_flag = pc_io_out_ex_io_br_io_br_flag; // @[Top.scala 57:29]
  assign if_io_reg_io_in_ex_io_br_io_br_target = pc_io_out_ex_io_br_io_br_target; // @[Top.scala 57:29]
  assign if_io_reg_io_stall_io_stall_flag = stall_io_out_stall_flag; // @[Top.scala 54:29]
  assign if_io_reg_io_stall_io_pred_miss_flag = stall_io_out_pred_miss_flag; // @[Top.scala 54:29]
  assign if_io_reg_n_clock = clock;
  assign if_io_reg_n_reset = reset;
  assign if_io_reg_n_io_in_reg_pc = if_io_reg_io_out_reg_pc; // @[Top.scala 45:29]
  assign if_io_reg_nn_clock = clock;
  assign if_io_reg_nn_reset = reset;
  assign if_io_reg_nn_io_in_reg_pc = if_io_reg_n_io_out_reg_pc; // @[Top.scala 67:29]
  assign id_io_reg_clock = clock;
  assign id_io_reg_reset = reset;
  assign id_io_reg_io_in_op1_data = id_io_out_op1_data; // @[Top.scala 63:25]
  assign id_io_reg_io_in_op2_data = id_io_out_op2_data; // @[Top.scala 63:25]
  assign id_io_reg_io_in_rd_addr = id_io_out_rd_addr; // @[Top.scala 63:25]
  assign id_io_reg_io_in_csr_addr_default = id_io_out_csr_addr_default; // @[Top.scala 63:25]
  assign id_io_reg_io_in_exe_fun = id_io_out_exe_fun; // @[Top.scala 63:25]
  assign id_io_reg_io_in_mem_wen = id_io_out_mem_wen; // @[Top.scala 63:25]
  assign id_io_reg_io_in_rd_wen = id_io_out_rd_wen; // @[Top.scala 63:25]
  assign id_io_reg_io_in_rd_sel = id_io_out_rd_sel; // @[Top.scala 63:25]
  assign id_io_reg_io_in_csr_cmd = id_io_out_csr_cmd; // @[Top.scala 63:25]
  assign id_io_reg_io_in_rs2_data = id_io_out_rs2_data; // @[Top.scala 63:25]
  assign id_io_reg_io_in_imm_b_sext = id_io_out_imm_b_sext; // @[Top.scala 63:25]
  assign id_io_reg_n_clock = clock;
  assign id_io_reg_n_reset = reset;
  assign id_io_reg_n_io_in_op1_data = id_io_reg_io_out_op1_data; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_op2_data = id_io_reg_io_out_op2_data; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_rd_addr = id_io_reg_io_out_rd_addr; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_csr_addr_default = id_io_reg_io_out_csr_addr_default; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_exe_fun = id_io_reg_io_out_exe_fun; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_mem_wen = id_io_reg_io_out_mem_wen; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_rd_wen = id_io_reg_io_out_rd_wen; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_rd_sel = id_io_reg_io_out_rd_sel; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_csr_cmd = id_io_reg_io_out_csr_cmd; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_rs2_data = id_io_reg_io_out_rs2_data; // @[Top.scala 69:29]
  assign id_io_reg_n_io_in_imm_b_sext = id_io_reg_io_out_imm_b_sext; // @[Top.scala 69:29]
  assign ex_io_reg_clock = clock;
  assign ex_io_reg_reset = reset;
  assign ex_io_reg_io_in_alu_io_alu_out = ex_io_out_alu_io_alu_out; // @[Top.scala 71:25]
  assign ex_io_reg_io_in_csr_io_csr_rdata = ex_io_out_csr_io_csr_rdata; // @[Top.scala 71:25]
  assign mem_io_reg_clock = clock;
  assign mem_io_reg_reset = reset;
  assign mem_io_reg_io_in_rd_wen = mem_io_out_rd_wen; // @[Top.scala 77:29]
  assign mem_io_reg_io_in_rd_addr = mem_io_out_rd_addr; // @[Top.scala 77:29]
  assign mem_io_reg_io_in_rd_data = mem_io_out_rd_data; // @[Top.scala 77:29]
endmodule
